library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package itc108_2_const is
	constant key_stop : integer := 1;
	constant key_rst : integer := 2;
	constant key_start : integer := 3;
	constant key_ok : integer := 5;
	constant key_down : integer := 6;
	constant key_up : integer := 7;
end package;
