-- graphics processing unit for the LCD display

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.itc.all;
use work.itc_lcd.all;

entity gpu is
	port (
		-- system
		clk   : in std_logic;
		rst_n : in std_logic;
		-- lcd
		l_addr : in l_addr_t;
		l_data : out l_px_t;
		-- program memory
		p_addr : out p_addr_t;
		p_data : in p_inst_t;
		-- image memory
		i_addr : out l_addr_t;
		i_data : in l_px_t; 
		-- user logic
		load  : in p_addr_t; -- load address in the program memory, value defined by constants generated by GIG
		ena  : in std_logic;
		busy : out std_logic
	);
end gpu;

architecture arch of gpu is

	signal start : std_logic;

	type state is (idle, foo);
begin

	edge_inst : entity work.edge(arch)
		port map(
			clk     => clk,
			rst_n   => rst_n,
			sig_in  => ena,
			rising  => start,
			falling => open
		);

	process (clk, rst_n) begin
		if rst_n = '0' then
			state <= idle;
		elsif rising_edge(clk) then
			case state is
				when idle =>
					if start = '1' then
						state <= foo;
					end if;
				when foo =>
					-- do something
				when others =>
					null;
			end case;
		end if;
	end process;

end arch;
