library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.itc.all;

package itc_lcd is
	constant lcd_width : integer := 128;
	constant lcd_height : integer := 160;
	constant lcd_color_depth : integer := 12;
	constant lcd_pixel_cnt : integer := lcd_width * lcd_height;
	constant lcd_bit_cnt : integer := lcd_pixel_cnt * lcd_color_depth;

	subtype pixel_t is unsigned(lcd_color_depth - 1 downto 0);
	type pixels_t is array (0 to lcd_pixel_cnt - 1) of pixel_t;

	--------------------------------------------------------------------------------
	-- command constants
	-- only the used commands are listed here
	--------------------------------------------------------------------------------

	constant lcd_slpout : u8_t := x"11";
	constant lcd_frmctr1 : u8_t := x"b1";
	constant lcd_pwctr1 : u8_t := x"c0";
	constant lcd_pwctr2 : u8_t := x"c1";
	constant lcd_pwctr3 : u8_t := x"c2";
	constant lcd_vmctr1 : u8_t := x"c5";
	constant lcd_gmctrp1 : u8_t := x"e0"; -- aka gamctrp1
	constant lcd_gmctrn1 : u8_t := x"e1"; -- aka gamctrn1
	constant lcd_colmod : u8_t := x"3a";
	constant lcd_dispon : u8_t := x"29";
	constant lcd_ramwr : u8_t := x"2c";

	--------------------------------------------------------------------------------
	-- initialization commands and arguments
	--------------------------------------------------------------------------------

	constant lcd_cmd_delay : u8_t := x"80";
	constant lcd_init : u8_arr_t(0 to 52) := (
		lcd_frmctr1, x"05", x"3c", x"3c",
		lcd_pwctr1, x"28", x"08", x"04",
		lcd_pwctr2, x"c0",
		lcd_pwctr3, x"0d", x"00",
		lcd_vmctr1, x"1a",
		lcd_gmctrp1, x"04", x"22", x"07", x"0a", x"2e", x"30", x"25", x"2a", x"28", x"26", x"2e", x"3a", x"00", x"01", x"03", x"13",
		lcd_gmctrn1, x"04", x"16", x"06", x"0d", x"2d", x"26", x"23", x"27", x"27", x"25", x"2d", x"3b", x"00", x"01", x"04", x"13",
		lcd_colmod, x"03",
		lcd_dispon,
		lcd_ramwr
	);
	constant lcd_init_dc : std_logic_vector(0 to 52) := not "10001000101001010000000000000000100000000000000001011";

	--------------------------------------------------------------------------------
	-- functions
	--------------------------------------------------------------------------------

	-- to_bytes: convert pixels_t to u8_arr_t
	-- pixels: array of pixels to convert
	function to_bytes(pixels : pixels_t) return u8_arr_t;

	--------------------------------------------------------------------------------
	-- font
	-- HD44780 5x7 pixel font data, http://eleif.net/HD44780.html 
	-- Array index is the relative ASCII code
	--------------------------------------------------------------------------------

	type glyph_t is array (0 to 6) of std_logic_vector(0 to 4);
	type font_t is array(32 to 127) of glyph_t;

	constant lcd_font : font_t := (-- this comment is for the formatter
	("00000", "00000", "00000", "00000", "00000", "00000", "00000"), -- [ 32] ' '
	("00100", "00100", "00100", "00100", "00000", "00000", "00100"), -- [ 33] '!'
	("01010", "01010", "01010", "00000", "00000", "00000", "00000"), -- [ 34] '"'
	("01010", "01010", "11111", "01010", "11111", "01010", "01010"), -- [ 35] '#'
	("00100", "01111", "10100", "01110", "00101", "11110", "00100"), -- [ 36] '
	("11000", "11001", "00010", "00100", "01000", "10011", "00011"), -- [ 37] '%'
	("01100", "10010", "10100", "01000", "10101", "10010", "01101"), -- [ 38] '&'
	("01100", "00100", "01000", "00000", "00000", "00000", "00000"), -- [ 39] '''
	("00010", "00100", "01000", "01000", "01000", "00100", "00010"), -- [ 40] '('
	("01000", "00100", "00010", "00010", "00010", "00100", "01000"), -- [ 41] ')'
	("00000", "00100", "10101", "01110", "10101", "00100", "00000"), -- [ 42] '*'
	("00000", "00100", "00100", "11111", "00100", "00100", "00000"), -- [ 43] '+'
	("00000", "00000", "00000", "00000", "01100", "00100", "01000"), -- [ 44] ','
	("00000", "00000", "00000", "11111", "00000", "00000", "00000"), -- [ 45] '-'
	("00000", "00000", "00000", "00000", "00000", "01100", "01100"), -- [ 46] '.'
	("00000", "00001", "00010", "00100", "01000", "10000", "00000"), -- [ 47] '/'
	("01110", "10001", "10011", "10101", "11001", "10001", "01110"), -- [ 48] '0'
	("00100", "01100", "00100", "00100", "00100", "00100", "01110"), -- [ 49] '1'
	("01110", "10001", "00001", "00010", "00100", "01000", "11111"), -- [ 50] '2'
	("11111", "00010", "00100", "00010", "00001", "10001", "01110"), -- [ 51] '3'
	("00010", "00110", "01010", "10010", "11111", "00010", "00010"), -- [ 52] '4'
	("11111", "10000", "11110", "00001", "00001", "10001", "01110"), -- [ 53] '5'
	("00110", "01000", "10000", "11110", "10001", "10001", "01110"), -- [ 54] '6'
	("11111", "10001", "00001", "00010", "00100", "00100", "00100"), -- [ 55] '7'
	("01110", "10001", "10001", "01110", "10001", "10001", "01110"), -- [ 56] '8'
	("01110", "10001", "10001", "01111", "00001", "00010", "01100"), -- [ 57] '9'
	("00000", "01100", "01100", "00000", "01100", "01100", "00000"), -- [ 58] ':'
	("00000", "01100", "01100", "00000", "01100", "00100", "01000"), -- [ 59] ';'
	("00010", "00100", "01000", "10000", "01000", "00100", "00010"), -- [ 60] '<'
	("00000", "00000", "11111", "00000", "11111", "00000", "00000"), -- [ 61] '='
	("01000", "00100", "00010", "00001", "00010", "00100", "01000"), -- [ 62] '>'
	("01110", "10001", "00001", "00010", "00100", "00000", "00100"), -- [ 63] '?'
	("01110", "10001", "00001", "01101", "10101", "10101", "01110"), -- [ 64] '@'
	("01110", "10001", "10001", "10001", "11111", "10001", "10001"), -- [ 65] 'A'
	("11110", "10001", "10001", "11110", "10001", "10001", "11110"), -- [ 66] 'B'
	("01110", "10001", "10000", "10000", "10000", "10001", "01110"), -- [ 67] 'C'
	("11100", "10010", "10001", "10001", "10001", "10010", "11100"), -- [ 68] 'D'
	("11111", "10000", "10000", "11110", "10000", "10000", "11111"), -- [ 69] 'E'
	("11111", "10000", "10000", "11110", "10000", "10000", "10000"), -- [ 70] 'F'
	("01110", "10001", "10000", "10111", "10001", "10001", "01111"), -- [ 71] 'G'
	("10001", "10001", "10001", "11111", "10001", "10001", "10001"), -- [ 72] 'H'
	("01110", "00100", "00100", "00100", "00100", "00100", "01110"), -- [ 73] 'I'
	("00111", "00010", "00010", "00010", "00010", "10010", "01100"), -- [ 74] 'J'
	("10001", "10010", "10100", "11000", "10100", "10010", "10001"), -- [ 75] 'K'
	("10000", "10000", "10000", "10000", "10000", "10000", "11111"), -- [ 76] 'L'
	("10001", "11011", "10101", "10101", "10001", "10001", "10001"), -- [ 77] 'M'
	("10001", "10001", "11001", "10101", "10011", "10001", "10001"), -- [ 78] 'N'
	("01110", "10001", "10001", "10001", "10001", "10001", "01110"), -- [ 79] 'O'
	("11110", "10001", "10001", "11110", "10000", "10000", "10000"), -- [ 80] 'P'
	("01110", "10001", "10001", "10001", "10101", "10010", "01101"), -- [ 81] 'Q'
	("11110", "10001", "10001", "11110", "10100", "10010", "10001"), -- [ 82] 'R'
	("01111", "10000", "10000", "01110", "00001", "00001", "11110"), -- [ 83] 'S'
	("11111", "00100", "00100", "00100", "00100", "00100", "00100"), -- [ 84] 'T'
	("10001", "10001", "10001", "10001", "10001", "10001", "01110"), -- [ 85] 'U'
	("10001", "10001", "10001", "10001", "10001", "01010", "00100"), -- [ 86] 'V'
	("10001", "10001", "10001", "10101", "10101", "10101", "01010"), -- [ 87] 'W'
	("10001", "10001", "01010", "00100", "01010", "10001", "10001"), -- [ 88] 'X'
	("10001", "10001", "10001", "01010", "00100", "00100", "00100"), -- [ 89] 'Y'
	("11111", "00001", "00010", "00100", "01000", "10000", "11111"), -- [ 90] 'Z'
	("11100", "10000", "10000", "10000", "10000", "10000", "11100"), -- [ 91] '['
	("10001", "01010", "11111", "00100", "11111", "00100", "00100"), -- [ 92] '\'
	("01110", "00010", "00010", "00010", "00010", "00010", "01110"), -- [ 93] ']'
	("00100", "01010", "10001", "00000", "00000", "00000", "00000"), -- [ 94] '^'
	("00000", "00000", "00000", "00000", "00000", "00000", "11111"), -- [ 95] '_'
	("01000", "00100", "00010", "00000", "00000", "00000", "00000"), -- [ 96] '`'
	("00000", "00000", "01110", "00001", "01111", "10001", "01111"), -- [ 97] 'a'
	("10000", "10000", "10110", "11001", "10001", "10001", "11110"), -- [ 98] 'b'
	("00000", "00000", "01110", "10000", "10000", "10001", "01110"), -- [ 99] 'c'
	("00001", "00001", "01101", "10011", "10001", "10001", "01111"), -- [100] 'd'
	("00000", "00000", "01110", "10001", "11111", "10000", "01110"), -- [101] 'e'
	("00110", "01001", "01000", "11100", "01000", "01000", "01000"), -- [102] 'f'
	("00000", "01111", "10001", "10001", "01111", "00001", "01110"), -- [103] 'g'
	("10000", "10000", "10110", "11001", "10001", "10001", "10001"), -- [104] 'h'
	("00100", "00000", "01100", "00100", "00100", "00100", "01110"), -- [105] 'i'
	("00010", "00000", "00110", "00010", "00010", "10010", "01100"), -- [106] 'j'
	("10000", "10000", "10010", "10100", "11000", "10100", "10010"), -- [107] 'k'
	("01100", "00100", "00100", "00100", "00100", "00100", "01110"), -- [108] 'l'
	("00000", "00000", "11010", "10101", "10101", "10001", "10001"), -- [109] 'm'
	("00000", "00000", "10110", "11001", "10001", "10001", "10001"), -- [110] 'n'
	("00000", "00000", "01110", "10001", "10001", "10001", "01110"), -- [111] 'o'
	("00000", "00000", "11110", "10001", "11110", "10000", "10000"), -- [112] 'p'
	("00000", "00000", "01101", "10011", "01111", "00001", "00001"), -- [113] 'q'
	("00000", "00000", "10110", "11001", "10000", "10000", "10000"), -- [114] 'r'
	("00000", "00000", "01110", "10000", "01110", "00001", "11110"), -- [115] 's'
	("01000", "01000", "11100", "01000", "01000", "01001", "00110"), -- [116] 't'
	("00000", "00000", "10001", "10001", "10001", "10011", "01101"), -- [117] 'u'
	("00000", "00000", "10001", "10001", "10001", "01010", "00100"), -- [118] 'v'
	("00000", "00000", "10001", "10101", "10101", "10101", "01010"), -- [119] 'w'
	("00000", "00000", "10001", "01010", "00100", "01010", "10001"), -- [120] 'x'
	("00000", "00000", "10001", "10001", "01111", "00001", "01110"), -- [121] 'y'
	("00000", "00000", "11111", "00010", "00100", "01000", "11111"), -- [122] 'z'
	("00010", "00100", "00100", "01000", "00100", "00100", "00010"), -- [123] '{'
	("00100", "00100", "00100", "00100", "00100", "00100", "00100"), -- [124] '|'
	("01000", "00100", "00100", "00010", "00100", "00100", "01000"), -- [125] '}'
	("00000", "00100", "00010", "11111", "00010", "00100", "00000"), -- [126] '~' -- right arrow
	("00000", "00100", "01000", "11111", "01000", "00100", "00000") --  [127] '' -- left arrow
	);
end package;

package body itc_lcd is
	function to_bytes(pixels : pixels_t) return u8_arr_t is
		variable joined_bits : unsigned(lcd_bit_cnt - 1 downto 0);
		variable result : u8_arr_t(lcd_bit_cnt / 8 - 1 downto 0);
	begin
		for p in pixels'range loop -- join into bits
			joined_bits(p * pixel_t'length + pixel_t'high downto p * pixel_t'length) := pixels(p);
		end loop;

		for b in result'range loop -- split info bytes
			result(b) := joined_bits(b * 8 + 7 downto b * 8);
		end loop;

		return result;
	end function;
end package body;
