--109工科技藝競賽數位電子職種
--術科參考試題一:裝置測試平台
--109.7.xx
--DHT11溫濕度感測器測試:1 wire
--TSL2561 I2C光感測器測試
--k4x4:
--0:啟動鍵, 1:重置鍵, 2:停止鍵, 4:上鍵, 5:下鍵, 6:確認鍵
--TFT_LCD128x160(132x162)(st7735)

--SD178BMI2C 語音播放模組
--SD178B address = 0b0100 000 (7 bits)
--SD178BMI2C指令表
--80H:停止、結束(即時執行命令碼)(V2版會死當)
--81H:增加音量0.5db(即時執行命令碼)
--82H:減少音量0.5db(即時執行命令碼)
--送完每個即刻執行的命令碼後，須等20ms後，才能再傳送I2C資料
--===========================================================
--以下2019 02 12 V2.2 版(修正舊版錯誤及新增指令)
--新增8F xx 2byte 指令
--02 8F 00 --Pause暫停
--02 8F 01 --Resume取消暫停
--02 8F 02 --Skip 提前結束正執行的87H或88H指令，跳至下一指令
--02 8F 03 --Soft Reset 重新開機
--
--===========================================================
--83H U8:調整播放速度比原始速度快U8%(00H~28H=0~40%)
--86H U8:設定輸出音量大小為U8(FFH FEH~01H 00H:0db,-0.5db,...,-127db,靜音無聲)預設音量值為D2H
--87H U32:延遲U32 ms時間(單位:ms)(高byte~低byte 00H00H00H80H=128ms)
--88H U16A U16B:播放microSD卡的wave音檔(U16A為檔名:1001~9999.wav 03E9H~270FH ,U16B:為循環播放次數，0表示無限次)
--1001:03E9,2000:07D0,3000:0BB8,4000:0FA0,5000:1388,6000:1770,7000:1B58,8000:1F40,9000:2328
--8AH U8:控制輸出接腳MO2~MO0狀態(U8[b2:b0]對應MO2~MO0狀態)

--8BH U8:Audio Amplifier WM8960 輸出通道控制
--	        WM8960 Audio 輸出通道開/關表
--通道	 Line Out 	  耳機		      喇叭
--代號	HP_R  HP_L 	HP_R  HP_L	 SPK_RN  SPK_LN
--U8	   AGND	 	OUT3(HP_C)	 SPK_RP  SPK_LP
--01H 	...................................Ⅴ
--02H 	...........................Ⅴ
--03H 	...........................Ⅴ......Ⅴ
--04H 	.............Ⅴ....Ⅴ
--05H 	...................Ⅴ..............Ⅴ
--06H 	.............Ⅴ............Ⅴ
--07H(預設)..........Ⅴ....Ⅴ......Ⅴ......Ⅴ
--08H 	.Ⅴ...Ⅴ
--09H 	......Ⅴ...........................Ⅴ
--0AH 	.Ⅴ........................Ⅴ
--0BH 	.Ⅴ...Ⅴ...................Ⅴ......Ⅴ

--109.7.xx版
--creator bye YHGL

--請使用秉華科技有限公司 TEL:04-26528352 www.be-friend.com.tw
--產品編號:BF-CYC3-S16A (EP3C16Q240C8 50MHz LEs:15,408 PINs:161)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

-- -----------------------------------------------------
entity E109_01_01 is
port(SCLK,S_RESET:in std_logic;			--系統 clk,reset

	 M7_0:in std_logic_vector(7 downto 0);--指撥開關 32xxxx10

	 --DHT11
	 DHT11_D_io:inout std_logic;		--DHT11 i/o

	 --LIGHT-TO-DIGITAL CONVERTER TSL2561
	 TSL2561_SCL:out std_logic;			--介面IO:SCL,如有接提升電阻時可設成inout
	 TSL2561_SDA:inout std_logic;		--介面IO:SDA,有接提升電阻
	 TSL2561_INT:in std_logic;			--TSL2561 INT

	 --k4x4鍵盤
	 ko:buffer std_logic_vector(3 downto 0);--偵測掃瞄線
	 ki:in std_logic_vector(3 downto 0);	--檢查回饋線
	 koo:buffer std_logic;					--觀察用(可有可無或不接線)

	 --D7S
	 SCANo:buffer std_logic_vector(7 downto 0);	--掃瞄信號
	 D7LED:out std_logic_vector(7 downto 0);	--顯示資料
     D7LED2:out std_logic_vector(7 downto 0);
     
	 --SD178BMI2C
	 SD178BMI2CP_3_3V_power:out std_logic_vector(7 downto 0);
	 SD178BMI2C_SCL:out std_logic;			--介面IO:SCL,如有接提升電阻時可設成inout
	 SD178BMI2C_SDA:inout std_logic;		--介面IO:SDA,有接提升電阻
	 SD178BMI2Co_reset:buffer std_logic:='1';--/reset
	 SD178BMI2Ci_MO0:in std_logic;			--/MO0

	 --tft_lcd_st7735_4w(CS,DC,SCL,SDA)+RES+BL----1.8'133x162 RGB TFT_LCD--108.07.20
     st7735_RESX:out std_logic;				--介面IO:RESx輸出
     st7735_CS:buffer std_logic;			--介面IO:CSx輸出
     st7735_DC:out std_logic;				--介面IO:DCx輸出
     st7735_SCL:buffer std_logic;			--介面IO:SCL輸出
     st7735_SDA:out std_logic;				--介面IO:SDA輸出
     st7735_BL:out std_logic;				--介面IO:SDA輸出

     --L293D DC motor 驅動IC
     --直流馬達可單向或雙向運轉驅動,或雙極性步進馬達驅動
     --輸出電流可達1A/L293 (600mA/L293D),電流要加倍時可將Y輸出並聯
     --目前使用方式:12組:直流馬達--34組:電源輸出控制(SD178BMI2C語音模組)
	 L293D_1A:buffer std_logic;		--介面IO:1A輸出:high ->1Y high
	 L293D_2A:buffer std_logic;		--介面IO:2A輸出:high ->2Y high
	 L293D_12EN:buffer std_logic;	--介面IO:12EN輸出:active high,low->1Y&2Y->Hz
	 L293D_3A:buffer std_logic;		--介面IO:3A輸出:high ->3Y high
	 L293D_4A:buffer std_logic;		--介面IO:4A輸出:high ->4Y high
	 L293D_34EN:buffer std_logic	--介面IO:34EN輸出:active high,low->3Y&4Y->Hz
    );
end E109_01_01;

-- -----------------------------------------------------
architecture YHGL of E109_01_01 is

	-- component=================================================================
	--tft_lcd_t7735 driver: 1.8'133x162 RGB TFT_LCD特急超飆速版
	component st7735_spi_tft_lcd_4w_driver_2 is
	   port(  st7735_CLK,st7735_RESET:in std_logic;		--系統時脈,系統重置
			  st7735_RES:in std_logic;					--介面控制:RESx輸入
			  st7735_BLS:in std_logic;					--介面控制:BL輸入
			  DCi:in std_logic_vector(1 downto 0);		--00:命令 01:命令參數 11:g資料
			  cmpai:in std_logic_vector(15 downto 0);	--命令_參數 輸入,水平16點image
			  cbi:in std_logic_vector(3 downto 0);		--色盤(4bit):xx01(12bit)、xx10(16bit)、xx11(18bit)
			  fcri,fcgi,fcbi:in std_logic_vector(7 downto 0);--色系
			  bcri,bcgi,bcbi:in std_logic_vector(7 downto 0);--色系
			  d8_1i:in integer range 0 to 16;			--水平剩餘點數1~16
			  --------------------------------------------------------------
			  st7735_RESX:out std_logic;				--介面IO:RESx輸出
			  st7735_CS:buffer std_logic;				--介面IO:CSx輸出
			  st7735_DC:out std_logic;					--介面IO:DCx輸出
			  st7735_SCL:buffer std_logic;				--介面IO:SCL輸出
			  st7735_SDA:out std_logic;					--介面IO:SDA輸出
			  st7735_BL:out std_logic;					--介面IO:BL輸出
			  --------------------------------------------------------------
			  st7735_reLOAD:out std_logic;				--載入旗標:0 可載入
			  st7735_LoadCK:in std_logic;				--載入時脈
			  st7735_spi_ok:buffer std_logic 			--完成旗標
			);
	end component st7735_spi_tft_lcd_4w_driver_2;
	signal st7735_CLK,st7735_RESET: std_logic;		--系統時脈,系統重置
	signal st7735_RES: std_logic;					--介面IO:RESx輸入
	signal st7735_BLS: std_logic;					--介面IO:BL輸入
	signal DCi: std_logic_vector(1 downto 0);		--00:命令 01:命令參數 11:g資料
	signal cmpai: std_logic_vector(15 downto 0);	--命令_參數 輸入,水平16點image
	signal cbi: std_logic_vector(3 downto 0);		--色盤(4bit):xx01(12bit)、xx10(16bit)、xx11(18bit)
	signal fcri,fcgi,fcbi: std_logic_vector(7 downto 0);--色系
	signal bcri,bcgi,bcbi: std_logic_vector(7 downto 0);--色系
	signal d8_1i:integer range 0 to 16;				--水平剩餘點數1~16
	signal st7735_reLOAD: std_logic;				--載入旗標:0 可載入
	signal st7735_LoadCK: std_logic;				--載入時脈
	signal st7735_spi_ok: std_logic;				--完成旗標

	---------------------------------------------------
	component k4x4 is
	port 
	(	kf,reset: in std_logic;
		ki: in std_logic_vector(3 downto 0);
		ko: buffer std_logic_vector(3 downto 0);
		kn,kv: buffer integer range 0 to 15;
		kok,koo: buffer std_logic	--koo測試觀察用169
	);
	end component;
	signal kf,kreset:std_logic;
	signal kn,kv:integer range 0 to 15;--鍵盤操作
	signal kok:std_logic;
	
	--DCmotor_pwm_driver=================================================================
	--pwmckset:設pwm範圍0~255,0:停止
	--pwmsetN:設pwm值 ,0:停止 ,0<pwmsetN>=pwmckset:100%全速運轉 ,1~pwmckset:pwm%
	--停止(0%):pwmckset=0
	--全速運轉(100%):pwmsetN>=pwmckset
	--pwm%=pwmsetN/pwmckset*100%
	--雙向運轉:?A?A輸入可控制停止(00,11)或正反轉(10,01),?EN可控制停止(0)或全速運轉或pwm%調速
	--單向運轉(原EN<-->A對調):?EN可控制停止(0)或運轉,?A?A輸入可控制停止(0)或全速運轉或pwm%調速
	component DCmotor_pwm_driver is
	port 
	(	DCmotor_CLK: in std_logic;					--驅動速率
		pwmckset,pwmsetN: in integer range 0 to 255;--pwmckset:設pwm範圍,pwmsetN:設pwm值
		A1,A2: in std_logic;						--轉向
		L293D_EN: out std_logic						--輸出
	);
	end component DCmotor_pwm_driver;
	signal pwmckset,pwmsetN:integer range 0 to 255;--pwmckset:設pwm範圍,pwmsetN:設pwm值
	constant DCmotor_base_pwm:integer range 0 to 63:=40;--最低轉速PWM設定值(1=0.5%pwm)

	--I2C_Driver--for TSL2561--------------------------------------------------------------
	component i2c2wdriver2
	Port(I2CCLK,RESET:in std_logic;					--系統時脈,系統重置
		ID:in std_logic_vector(3 downto 0);			--裝置碼
		CurrentADDR:in std_logic;					--要求命令:(0目前位址讀取),(1指定位址讀取)
		ADDR:in std_logic_vector(7 downto 0);		--位置(COMMAND)
		A2A1A0:in std_logic_vector(2 downto 0);		--位置,最多8個位址並存
		DATAin:in std_logic_vector(7 downto 0);		--資料輸入
		DATAout:buffer std_logic_vector(7 downto 0);--資料輸出
		RW:in std_logic;							--讀寫
		RWN:in integer range 0 to 15;				--嘗試讀寫次數
		D_W_R_N:in integer range 0 to 63;		 	--連續讀寫次數
		D_W_R_Nok:buffer std_logic;					--讀寫1次數旗標
		reWR:in std_logic;							--已寫入或讀出資料
		I2Cok,I2CS:buffer std_logic;				--I2Cok,CS 狀態
		SCL:out std_logic;							--介面IO:SCL,如有接提升電阻時可設成inout
		SDA:inout std_logic							--介面IO:SDA
		);
	end component;

	--TSL2561
	signal TSL2561_ID:std_logic_vector(3 downto 0):="0111";--TSL2561 ADDR SEL :(Float:0111,GND:0101,VDD:1001),24LCxx裝置碼:"1010"
	signal TSL2561_DATAin,TSL2561_DATAout:std_logic_vector(7 downto 0);
			--I2C時脈	,	啟動 	,I2C完成	,狀態		,讀寫
	signal TSL2561_CLK,TSL2561_RESET,TSL2561_ok,TSL2561_CS,TSL2561_RW:std_logic;--
	constant TSL2561_RWN:integer range 0 to 15 :=3;		--嘗試讀寫1次設定
	signal TSL2561_COMMAND:std_logic_vector(7 Downto 0);--位址(ADDR:COMMAND)
	signal TSL2561_D_W_R_N:integer range 0 to 63;		--page 長度
	signal TSL2561_reWR,TSL2561_D_W_R_Nok:std_logic;	--繼續,通知處理

	--------------------------------------------------------------------------------------	
	--DHT11_driver
	--Data format:
	--DHT11_DBo(std_logic_vector:8bit):由DHT11_RDp選取輸出項
	--RDp=5:chK_SUM
	--RDp=4							   3							   2								1								  0					
	--The 8bit humidity integer data + 8bit the Humidity decimal data +8 bit temperature integer data + 8bit fractional temperature data +8 bit parity bit.
	--直接輸出濕度(DHT11_DBoH)及溫度(DHT11_DBoT):integer(0~255:8bit),直接輸出溫度小數(DHT11_DBoT_1)
	--AOSONG版:起動較快速
	--(規格測試範圍:0~50℃、20~90%RH)無小數部分(全為0)
	--ASAIR版:起動較慢，所以須將驅動硬體有兩處做修改:11改為14即可
	--(規格測試範圍:-20~60℃ ?溫度小數部分第7位元表示0正1負、第3..0位元為0~9小數部分?、5~95%RH無小數部分)
	--可由DHT11_RDp=1 ->DHT11_DBo(溫度小數一位):DHT11_DBo(7)='1'->-T,DHT11_DBo(7)='0'->+T,DHT11_DBo(3 downto 0)=小數位數0~9

	component DHT11_driver is
		port
		(	DHT11_CLK,DHT11_RESET:in std_logic;		--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))操作速率,重置
			DHT11_D_io:inout std_logic;				--DHT11 i/o
			DHT11_DBo:out std_logic_vector(7 downto 0);--DHT11_driver 資料輸出
			DHT11_RDp:in integer range 0 to 7;		--資料讀取指標
			DHT11_tryN:in integer range 0 to 7;		--錯誤後嘗試幾次
			DHT11_ok,DHT11_S:buffer std_logic;		--DHT11_driver完成作業旗標,錯誤信息
			DHT11_DBoH,DHT11_DBoT,DHT11_DBoT_1:buffer integer range 0 to 255;--直接輸出濕度(整數,小數固定為0值所以不輸出),溫度(整數),溫度小數1位(bit7=1為負值)
			DHT11_DBoH1,DHT11_DBoH0,DHT11_DBoT1,DHT11_DBoT0,DHT11_DBoT_1_1:buffer integer range 0 to 9;--直接輸出濕度及溫度(十位數及個位數)
			DHT11_DBoH1_ASC,DHT11_DBoH0_ASC,DHT11_DBoT1_ASC,DHT11_DBoT0_ASC,DHT11_DBoT_1_1_ASC:buffer std_logic_vector(7 downto 0);--直接輸出濕度及溫度ASCII
			H_Sound_DATA,T_Sound_DATA:buffer std_logic_vector(31 downto 0)--直接輸出濕度及溫度語音
		);
	end component DHT11_driver;
	Signal DHT11_CLK,DHT11_RESET:std_logic;		--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))操作速率,重置
	Signal DHT11_DBo:std_logic_vector(7 downto 0);--DHT11_driver 資料輸出
	Signal DHT11_RDp:integer range 0 to 7:=1;	--資料讀取指標5~0,1:(溫度小數一位)
	Signal DHT11_tryN:integer range 0 to 7:=3;	--錯誤後嘗試幾次
	Signal DHT11_ok,DHT11_S:std_logic;			--DHT11_driver完成作業旗標,錯誤信息	
	Signal DHT11_DBoH,DHT11_DBoT,DHT11_DBoT_1:integer range 0 to 255;
	Signal DHT11_DBoH1,DHT11_DBoH0,DHT11_DBoT1,DHT11_DBoT0,DHT11_DBoT_1_1:integer range 0 to 9;
	Signal DHT11_DBoH1_ASC,DHT11_DBoH0_ASC,DHT11_DBoT1_ASC,DHT11_DBoT0_ASC,DHT11_DBoT_1_1_ASC:std_logic_vector(7 downto 0);
	Signal H_Sound_DATA,T_Sound_DATA:std_logic_vector(31 downto 0);--濕度及溫度語音

	-------------------------------------------------------------------------------------
	component sd178BMI2C2wdriver
	 port(I2CCLK,RESET:in std_logic;				--系統時脈,系統重置
		  ID:in std_logic_vector(6 downto 0);		--裝置碼0100000
		  DATAin:in std_logic_vector(7 downto 0);	--資料輸入
		  DATAout:buffer std_logic_vector(7 downto 0);--資料輸出
		  RW:in std_logic;							--讀寫
		  RWN:in integer range 0 to 15;				--嘗試讀寫次數
		  D_W_R_N:in integer range 0 to 255;	 	--連續讀寫次數
		  D_W_R_Nok:buffer std_logic;				--讀寫1次數旗標
		  reWR:in std_logic;						--已寫入或讀出資料
		  I2Cok,I2CS:buffer std_logic;				--I2Cok,CS 狀態
		  SCL:out std_logic;						--介面IO:SCL,如有接提升電阻時可設成inout
		  SDA:inout std_logic						--介面IO:SDA
		 );
	end component;
	--單筆操作:D_W_R_N=1
	--多筆操作:由D_W_R_N指定,每完成1筆回D_W_R_Nok,收到reWR後再進行下一筆

	--SD178BMI2C
	signal SD178BMI2C_ID:std_logic_vector(6 downto 0):="0100000";
	signal SD178BMI2C_DATAin,SD178BMI2C_DATAout:std_logic_vector(7 downto 0);
			--I2C時脈,			啟動		,I2C完成	,狀態			,讀寫
	signal SD178BMI2C_CLK,SD178BMI2C_RESET,SD178BMI2C_ok,SD178BMI2C_CS,SD178BMI2C_RW:std_logic;--
	constant SD178BMI2C_RWN:integer range 0 to 15 :=1;		--嘗試讀寫1次設定
	signal SD178BMI2C_D_W_R_N:integer range 0 to 255;		--page 長度
	signal SD178BMI2C_reWR,SD178BMI2C_D_W_R_Nok:std_logic;	--繼續,通知處理

	-------------------------------------------------------------------------------------
	type D7_T is array (7 downto 0) of integer range 0 to 17;
	signal D7_DB:D7_T;		--顯示資料
	signal d7dot,flashs,flash_a_g:std_logic_vector(7 downto 0);
	signal flash_a_gs:std_logic_vector(6 downto 0);
	signal scanP:integer range 0 to 7;	--掃瞄指標
	--BCD碼解共陽極七段顯示碼gfedcba
	type D7LED_T is array (0 to 16) of std_logic_vector(6 Downto 0);
	constant Disp7:D7LED_T:=("0111111",
							"0000110",
							"1011011",
							"1001111",
							"1100110",
							"1101101",
							"1111101",
							"0000111",
							"1111111",
							"1101111",
							"1111001",
							"1110001",
							"1110110",
							"0111000",
							"1110111",
							"0111110",
							"0000000");--16不顯示

	--TSL2561-----------------------------------------------------------------------------
	signal TSL2561P_reset,TSL2561P_ok:std_logic;
	signal TSL2561_DP:integer range 0 to 3;
	type TSL2561_DATA01_T is array (0 to 3) of std_logic_vector(7 downto 0);
	signal TSL2561_DATA01:TSL2561_DATA01_T;
	signal CH0,CH1:integer range 0 to 65535;
	signal Tint:integer range 0 to 3:=2;
	signal iGain,iType:integer range 0 to 1:=0;
	signal chScale0:std_logic_vector(15 downto 0);	--16bit
	signal chScale1:std_logic_vector(19 downto 0);	--20bit
	signal chScale:integer range 0 to 1048575;		--20bit 2^20-1
	type chScale_T is array (0 to 2) of std_logic_vector(15 downto 0);
	constant chScale_TS:chScale_T:=(X"7517",X"0FE7",X"0400");
	signal channe0:integer range 0 to 67108863;		--26bit 2^26-1
	signal channe1:std_logic_vector(25 downto 0);	--26bit
	signal ratio1:integer range 0 to 4095;			--12bit 2^12-1
	signal ratio:std_logic_vector(11 downto 0);		--12bit
	signal BM:integer range 0 to 7;
	type KTC_T is array (0 to 7) of std_logic_vector(11 downto 0);
	constant KT_T_FN_CL:KTC_T:=(X"040",X"080",X"0c0",X"100",X"138",X"19a",X"29a",X"29a");
	constant BT_T_FN_CL:KTC_T:=(X"1f2",X"214",X"23f",X"270",X"16f",X"0d2",X"018",X"000");
	constant MT_T_FN_CL:KTC_T:=(X"1be",X"2d1",X"37b",X"3fe",X"1fc",X"0fb",X"012",X"000");
	constant KT_CS:KTC_T:=(X"043",X"085",X"0c8",X"10a",X"14d",X"19a",X"29a",X"29a");
	constant BT_CS:KTC_T:=(X"204",X"228",X"253",X"282",X"177",X"101",X"037",X"000");
	constant MT_CS:KTC_T:=(X"1ad",X"2c1",X"363",X"3df",X"1dd",X"127",X"02b",X"000");
	signal KTC,BTC,MTC:KTC_T;
	signal tempb,tempm,temp0,temp:integer range 0 to 520093695;		--32bit :0~2^32-1
	signal LUXS,LUXS1,LUXS2,LUXS3:integer range 0 to 65535;	--16bit:0~2^16-1
	signal LUXSx,LUXSx1,LUXSx2:integer range 0 to 65535;	--16bit:0~2^16-1
	type LUX_T is array (0 to 3) of integer range 0 to 15;
	signal LUX:D7_T:=(0,0,0,0,0,0,0,0);	--顯示資料
	signal LUXDP:integer range 0 to 7;	--小數點位置

	-- tft lcd_st7735------------------------------------------------------------------------
	--st7735指令表格式:
	type st7735_T is array (0 to 27) of std_logic_vector(7 Downto 0);
	signal st7735_IT:st7735_T:=(X"11",	--0 Default SLPIN(10h), SLPOUT(11h), 120ms:--休眠/喚醒

								X"29", 	--1 DISPON (29h), Default DISPOFF (28h), 120ms:--顯示on/off

								X"B4", 	--2 INVCTR (B4h): Display Inversion Control:--反相控制
								X"03",  --3 Default(03h): 0 0 0 0 0 NLA NLB NLC: 00000011

								X"36", 	--4 MADCTL (36h): Memory Data Access Control:--記憶體進出入順序及顯示控制
								X"C0", 	--5 Default(00h): MY(0) MX(0) MV(0) ML(0) RGB(0) MH(0) - -

								X"38",	--6 Default IDMOFF (38h)(4k,65k,262k), IDMON (39h)(only 8 color):--色彩限定

								X"20", 	--7 Default INVOFF (20h): Display Inversion Off, INVON (21h): Display Inversion On:--不反相／反相顯示

								X"13",	--8 Default NORON (13h): Normal Display Mode On, PTLON (12h): Partial Display Mode On:--正常／部分顯示模式

								X"30", 	--9 PTLAR (30h): Partial Area:--顯示部分範圍設定
								X"00",	--10 PSL
								X"00",	--11
								X"00",	--12 PEL
								X"A1",	--13

								X"3A",	--14 COLMOD (3Ah): Interface Pixel Format:--色彩深度設定(12-bit,16-bit,18-bit)
								X"06",	--15 Default(06h):18 bit pixel format, (05h):16 bit pixel format, (03h):12 bit pixel format

								X"2A", 	--16 CASET (2Ah): Column Address Set, Default 0~131:132:--frame x範圍設定0~131共132
								X"00",  --17 XS
								X"00",  --18
								X"00", 	--19 XE
								X"83",  --20 (131)

								X"2B", 	--21 RASET (2Bh): Row Address Set, Default 0~161:162:--frame y範圍設定0~161共162
								X"00",  --22 YS
								X"00",  --23
								X"00",  --24 YE
								X"A1",  --25 (161)

								X"2C", 	--26 RAMWR (2Ch): Memory Write:--寫入顯示資料
								
								X"28" 	--27 user defined region(must expand on its own):DISPON (29h), Default DISPOFF (28h), 120ms:--顯示on/off,
								);

	type st7735_cT0 is array (0 to 2) of std_logic_vector(7 Downto 0);--(R,G,B)
	type st7735_cT1 is array (0 to 9) of st7735_cT0;
	signal st7735_8baseCOLOR:st7735_cT1:=((X"00",X"00",X"00"),--0 BLACK
										  (X"FF",X"00",X"00"),--1 RED
										  (X"00",X"FF",X"00"),--2 GREEN
										  (X"00",X"00",X"FF"),--3 BLUE
										  (X"FF",X"FF",X"00"),--4 YELLOW
										  (X"FF",X"00",X"FF"),--5 MAGENTA
										  (X"00",X"FF",X"FF"),--6 CYAN
										  (X"FF",X"FF",X"FF"),--7 WHITE
										  (X"00",X"00",X"00"),--8 user defined
										  (X"00",X"00",X"00"));--9user defined

	signal B1_COLORi,B0_COLORi,monoC:integer range 0 to 9;

	signal st7735_DATA_C_INC:integer range 0 to 16;
	signal st7735_COM_PN,st7735_COM_PN0:integer range 0 to 31;
	signal st7735_COM_POINTER,st7735_COM_POINTERs:integer range 0 to 127;
	signal st7735_P_CLK,st7735_P_RESET,st7735_P_ok:std_logic;
	signal st7735_reset0:std_logic;--啟動TFT_LCD首次清空
	
	signal gdata,gdata0,gdata1,gdata2,gdata3,gdata4,gdata5,gdata6,gdata7:std_logic_vector(15 Downto 0);
	signal gdata8,gdata9,gdata10,gdata11,gdata12,gdata13,gdata14,gdata15:std_logic_vector(15 Downto 0);
	signal fc2,bc2:st7735_cT0:=(X"00",X"00",X"00");
	signal cbis:std_logic_vector(3 Downto 0);
	signal st7735_ch:std_logic_vector(3 Downto 0);	
	
	signal st7735_COLMOD,st7735_INVCTR,st7735_MADCTL,st7735_IDMOFF_ON:std_logic_vector(7 Downto 0);
	signal st7735_INVOFF_ON,st7735_NORON_PTLON,st7735_DISPON_OFF:std_logic_vector(7 Downto 0);
	signal st7735_PSL,st7735_PEL:integer range 0 to 255;
	signal st7735_DATA_CPOINTER,st7735_DATA_RPOINTER:integer range 0 to 255;
	signal st7735_DATA_CPOINTER_begin,st7735_DATA_CPOINTER_end,st7735_x,st7735_xincN:integer range 0 to 255;
	signal st7735_DATA_RPOINTER_begin,st7735_DATA_RPOINTER_end,st7735_y:integer range 0 to 255;
	signal st7735_xinc1:integer range 0 to 32767;
	signal st7735_time_Dn:integer range 0 to 100000000;--2s
	signal isword:boolean:=false;				--圖形或字型?圖形
	signal word_w,W_w_b:integer range 0 to 127;	--字寬,bit餘數
	signal st7735_x0:integer range 0 to 3;		--去前導零xxx.x
	signal remove_leading_0:std_logic;			--去前導零on/off
	type st7735_DATA_T is array (0 to 4) of integer range 0 to 9;
	signal st7735_DATA:st7735_DATA_T;

	-- -----------------------------------------------------
	--SD178BMI2C			 設語音表長度
	type SD178BMI2C_T is array (0 to 255) of std_logic_vector(7 downto 0);
	signal SD178BMI2C_sound:SD178BMI2C_T;			--(0:語音播放長度),....
	signal SD178BMI2CP_reseton_delay:integer range 0 to 255;--power on delay
	signal SD178BMI2C_IL:integer range 0 to 255;	--語音表取值指標
	signal SD178BMI2CP_reset,SD178BMI2CP_ok,SD178BMI2C_RWs:std_logic;--SD178BMI2CP 重置 ,完成 ,讀寫(1:read,0:write)
	signal SD178BMI2CP_powerdown,SD178BMI2CP_reseton:std_logic;--power on/off,RESET
	signal SD178BMI2C_P_end_t_onoff:std_logic:='0';				--是否啟動終止延遲計時
	signal SD178BMI2C_P_end_t_set:integer range 0 to 32767:=0;	--終止延遲計時次數(1:約1.004ms)
	type SD178BMI2C_rT is array (0 to 4) of std_logic_vector(7 downto 0);
	signal SD178BMI2C_DATA0_4:SD178BMI2C_rT;

	signal Sound88:std_logic_vector(7 downto 0);
	constant Soundclr80:std_logic_vector(7 downto 0):=X"80";	--清除SD178B buffer內的所有碼,停止正在執行的動作,已執行的設定不變(2.0V會當機)
	constant Soundup81:std_logic_vector(7 downto 0):=X"81";		--音量遞增即時指令
	constant Sounddown82:std_logic_vector(7 downto 0):=X"82";	--音量遞減即時指令
	--音量表
	type Sound86_90_VOT is array (0 to 9) of std_logic_vector(7 downto 0);
	--constant Sound86_90:Sound86_90_VOT:=(X"00",X"87",X"96",X"A5",X"B4",X"C3",X"D2",X"E1",X"F0",X"FF");--音量表
	constant Sound86_VOL:Sound86_90_VOT:=(X"00",X"C0",X"C8",X"D0",X"D8",X"E0",X"E8",X"F0",X"F8",X"FF");--音量表
	--聲道表
	--HP_R-HP_L		:100-LR:靠靜音關閉 :101-L,110-R,111-LR
	--SPK_RN-SPK_LN :100-xx(可以全關掉):101-L,110-R,111-LR
	type Sound8B_R_L_T is array (0 to 3) of std_logic_vector(7 downto 0);
	constant Sound8B_R_L:Sound8B_R_L_T:=(X"04",X"06",X"05",X"07");--聲道表
	
	signal F12:integer range 0 to 1;--01功能選項
	signal F1,Sound86:integer range 0 to 9;--音量選項
	signal F2,Sound8B:integer range 0 to 3;--聲道選項

	-- -----------------------------------------------------
	signal FD:std_logic_vector(25 downto 0);					 --除頻器
	signal SW_CLK,E109_1_1_MainCLK,OLED_P_CLK,OLED_P_RESET:std_logic;--防彈跳時脈,主控器操控頻率,OLED
	--計時計數
	signal times:integer range 0 to 4095;
	signal times1:integer range 0 to 511;
	signal S0on:std_logic;
	--指撥開關
	type M7_0T is array (0 to 7) of std_logic_vector(2 downto 0);
	signal M70s:M7_0T;
	signal M710,MMx,MM:std_logic_vector(1 downto 0);
	signal M776:std_logic_vector(1 downto 0);
	signal MMs,soundn:integer range 0 to 7;
	signal Mx:std_logic_vector(3 downto 0);

	--==tft lcd 圖形===================================================================================
	--字型&圖形 16bit
	signal beFriendC_P:integer range 0 to 16383;
	type beFriendt is array (0 to 16383) of integer range 0 to 65535;--(0,2^14-1)16bit
	constant beFriend:beFriendt:=
	(
	--20x40字:2x40=80
	--0:0:79
	0,0,0,0,0,0,0,0,0,0,1016,0,3900,0,7710,0,7695,0,15367,32768,15367,32768,30727,32768,30723,49152,30723,49152,30723,49152,61443,49152,61443,49152,61443,49152,61443,57344,61443,57344,61443,57344,61443,57344,61443,49152,61443,49152,61443,49152,30723,49152,30723,49152,30723,49152,30727,32768,15367,32768,15367,0,7695,0,3614,0,1980,0,1008,0,0,0,0,0,0,0,0,0,0,0,
	--1:80:159
	0,0,0,0,0,0,0,0,0,0,48,0,240,0,1008,0,4080,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,112,0,120,0,248,0,2047,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--2:160:239
	0,0,0,0,0,0,0,0,0,0,1008,0,4092,0,7294,0,14399,0,12319,0,28687,0,28687,32768,24583,32768,57351,32768,7,32768,7,0,15,0,15,0,15,0,30,0,30,0,60,0,56,0,112,0,240,0,480,0,448,0,896,0,1792,0,3584,57344,7681,49152,7171,49152,16383,32768,65535,32768,0,0,0,0,0,0,0,0,0,0,0,0,
	--3:240:319
	0,0,0,0,0,0,0,0,0,0,1020,0,2046,0,3615,0,7183,0,7175,0,14343,32768,12295,32768,7,0,7,0,14,0,14,0,28,0,124,0,510,0,1023,0,15,32768,7,32768,3,49152,3,49152,3,49152,3,49152,1,49152,1,49152,3,32768,3,32768,7,0,15,0,15902,0,16376,0,8160,0,0,0,0,0,0,0,0,0,0,0,
	--4:320:399
	0,0,0,0,0,0,0,0,0,0,6,0,14,0,30,0,30,0,62,0,62,0,126,0,238,0,238,0,462,0,974,0,910,0,1806,0,1806,0,3598,0,7694,0,7182,0,14350,0,14350,0,28686,0,32767,57344,32767,57344,14,0,14,0,14,0,14,0,14,0,14,0,14,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--5:400:479
	0,0,0,0,0,0,0,0,0,49152,3,49152,1023,32768,1023,32768,896,0,1792,0,1792,0,3840,0,3584,0,3968,0,8176,0,8184,0,5118,0,126,0,31,0,15,32768,7,32768,7,32768,3,32768,3,49152,3,49152,3,49152,3,32768,3,32768,3,32768,7,0,7,0,14,0,32284,0,16376,0,8128,0,0,0,0,0,0,0,0,0,0,0,
	--6:480:559
	0,0,0,0,0,0,0,0,0,0,31,49152,124,0,240,0,992,0,1984,0,1920,0,3840,0,7680,0,7680,0,15360,0,15360,0,32766,0,32703,0,31759,32768,30727,32768,30727,49152,30723,49152,28675,49152,28675,49152,28675,49152,28675,49152,30723,49152,30723,49152,30723,49152,14339,49152,15363,32768,7687,32768,3855,0,2046,0,1016,0,0,0,0,0,0,0,0,0,0,0,
	--7:560:639
	0,0,0,0,0,0,0,0,0,0,8191,57344,16383,49152,14337,49152,14339,49152,28675,32768,24579,32768,7,32768,7,0,7,0,7,0,15,0,14,0,14,0,30,0,28,0,28,0,60,0,60,0,56,0,56,0,120,0,112,0,112,0,240,0,240,0,224,0,480,0,480,0,448,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--8:640:719
	0,0,0,0,0,0,0,0,0,0,508,0,1935,0,3591,32768,7171,32768,7171,49152,7171,49152,7171,49152,7171,49152,7683,32768,7687,32768,3847,0,3982,0,2044,0,1016,0,508,0,510,0,1983,0,3855,32768,3591,32768,7171,49152,7171,49152,15361,49152,15361,49152,15361,49152,15361,49152,7169,49152,7681,49152,3843,32768,1999,0,508,0,0,0,0,0,0,0,0,0,0,0,
	--9:720:799
	0,0,0,0,0,0,0,0,0,0,1016,0,1822,0,3599,0,7175,32768,7175,32768,15363,49152,14339,49152,14339,49152,30721,57344,30721,57344,30721,57344,30721,57344,31745,57344,15361,57344,15361,57344,7683,57344,7943,49152,4095,49152,1011,49152,3,49152,7,32768,7,32768,15,0,31,0,30,0,60,0,120,0,496,0,1984,0,16128,0,0,0,0,0,0,0,0,0,0,0,
	--.:800:879
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,240,0,504,0,504,0,504,0,240,0,0,0,0,0,0,0,0,0,0,0,
	--32x40:2x40=80
	--space: 880:959
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--O:960:1039
	0,0,0,0,0,0,0,0,0,0,31,61440,120,31744,240,7680,480,3840,960,1920,1920,960,3840,480,3840,480,7936,496,7680,240,7680,240,7680,240,7680,240,7680,240,15872,240,15872,248,7680,240,7680,240,7680,240,7680,240,7680,240,3840,480,3840,480,3968,992,1920,960,960,1920,480,3840,240,7680,124,31744,15,57344,0,0,0,0,0,0,0,0,0,0,
	--F:1040:1119
	0,0,0,0,0,0,0,0,0,0,0,0,2047,65472,248,960,240,448,240,448,240,192,240,64,240,0,240,0,240,1792,240,1792,240,1792,240,3840,240,7936,255,65280,240,3840,240,1792,240,1792,240,1792,240,0,240,0,240,0,240,0,240,0,240,0,240,0,248,0,248,0,2047,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--28x40:80
	--LUX.:1120:1199
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,28910,60928,8260,17408,8260,10240,8260,10240,8260,4096,8260,10240,8772,10240,9284,17408,31800,60992,0,0,0,0,0,0,0,0,0,0,0,0,
	--oC:1200:1279
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8064,0,14720,0,12736,49152,12751,65280,14748,3840,7992,1792,120,768,112,384,112,0,224,0,224,0,224,0,224,0,224,0,224,0,224,0,240,0,112,384,112,384,56,768,60,1792,30,3584,7,64512,0,0,0,0,0,0,0,0,0,0,
	--%:1280:1359
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,240,12288,508,61440,927,57344,1948,57344,1820,49152,3865,49152,3609,32768,3611,32768,3635,0,3703,0,2022,32512,974,62208,13,58112,29,49920,25,49920,59,50944,51,34304,115,34304,97,52224,225,55296,224,61440,0,0,0,0,0,0,0,0,0,0,
	
	--大字:123456789: 128/16*160=1280=1280*16bit=20480bit
	--1:1360:2639
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,768,0,0,0,0,0,0,0,3840,0,0,0,0,0,0,0,16128,0,0,0,0,0,0,0,65280,0,0,0,0,0,0,7,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,511,65280,0,0,0,0,0,0,4095,65280,0,0,0,0,0,0,16383,65280,0,0,0,0,0,0,65535,65280,0,0,0,
	0,0,3,65535,65280,0,0,0,0,0,31,65535,65280,0,0,0,0,0,127,65535,65280,0,0,0,0,0,511,65535,65280,0,0,0,0,0,2047,65535,65280,0,0,0,0,0,8191,65535,65280,0,0,0,0,0,8191,65535,65280,0,0,0,0,0,8191,65535,65280,0,0,0,0,0,8190,1023,65280,0,0,0,0,0,8128,511,65280,0,0,0,0,0,7168,255,65280,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,
	0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,255,65408,0,0,0,0,0,0,255,65408,0,0,0,0,0,0,255,65408,0,0,0,0,0,0,511,65408,0,0,0,0,0,0,511,65472,0,0,0,0,0,0,1023,65504,0,0,0,0,0,0,2047,65520,0,0,0,
	0,0,0,8191,65528,0,0,0,0,0,0,65535,65535,0,0,0,0,0,31,65535,65535,64512,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,2047,65535,65535,65528,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--2:2640:3919
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,127,61440,0,0,0,0,0,0,4095,65280,0,0,0,0,0,0,32767,65504,0,0,0,0,0,1,65535,65528,0,0,0,0,0,7,65535,65534,0,0,0,0,0,31,65535,65535,32768,0,0,0,0,127,65535,65535,49152,0,0,0,0,255,65535,65535,57344,0,0,0,0,511,65535,65535,61440,0,0,0,0,2047,65535,65535,64512,0,0,0,0,4095,65535,65535,65024,0,0,0,0,8191,65535,65535,65024,0,0,
	0,0,16383,65535,65535,65280,0,0,0,0,16383,65535,65535,65408,0,0,0,0,32767,61695,65535,65472,0,0,0,0,65535,3,65535,65504,0,0,0,1,65528,0,32767,65504,0,0,0,1,65520,0,8191,65520,0,0,0,3,65504,0,2047,65528,0,0,0,7,65408,0,1023,65528,0,0,0,7,65280,0,511,65532,0,0,0,15,65280,0,255,65532,0,0,0,15,65024,0,127,65534,0,0,0,31,64512,0,63,65534,0,0,0,31,63488,0,31,65535,0,0,0,63,63488,0,15,65535,0,0,0,63,61440,0,7,65535,0,0,0,63,61440,0,7,65535,32768,0,
	0,127,57344,0,3,65535,32768,0,0,127,57344,0,3,65535,32768,0,0,127,57344,0,1,65535,32768,0,0,255,49152,0,0,65535,49152,0,0,255,49152,0,0,65535,49152,0,0,255,32768,0,0,65535,49152,0,0,511,32768,0,0,32767,49152,0,0,511,0,0,0,32767,49152,0,0,511,0,0,0,16383,49152,0,0,511,0,0,0,16383,49152,0,0,1022,0,0,0,16383,49152,0,0,1022,0,0,0,16383,49152,0,0,1020,0,0,0,16383,49152,0,0,1020,0,0,0,8191,49152,0,0,2044,0,0,0,8191,49152,0,0,2040,0,0,0,8191,49152,0,
	0,2040,0,0,0,8191,49152,0,0,2040,0,0,0,8191,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,16383,49152,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,32767,0,0,0,0,0,0,0,32767,0,0,0,0,0,0,0,32767,0,0,
	0,0,0,0,0,32767,0,0,0,0,0,0,0,65535,0,0,0,0,0,0,0,65534,0,0,0,0,0,0,0,65534,0,0,0,0,0,0,1,65534,0,0,0,0,0,0,1,65532,0,0,0,0,0,0,3,65532,0,0,0,0,0,0,3,65532,0,0,0,0,0,0,3,65528,0,0,0,0,0,0,7,65528,0,0,0,0,0,0,7,65520,0,0,0,0,0,0,15,65520,0,0,0,0,0,0,15,65504,0,0,0,0,0,0,15,65504,0,0,0,0,0,0,31,65504,0,0,0,0,0,0,31,65472,0,0,
	0,0,0,0,63,65408,0,0,0,0,0,0,127,65408,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,255,65024,0,0,0,0,0,0,511,65024,0,0,0,0,0,0,511,64512,0,0,0,0,0,0,1023,63488,0,0,0,0,0,0,2047,63488,0,0,0,0,0,0,2047,61440,0,0,0,0,0,0,4095,61440,0,0,0,0,0,0,4095,57344,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,16383,32768,0,0,0,0,0,0,32767,0,0,0,
	0,0,0,0,65534,0,0,0,0,0,0,1,65532,0,0,0,0,0,0,1,65532,0,0,0,0,0,0,3,65528,0,0,0,0,0,0,7,65520,0,0,0,0,0,0,7,65504,0,0,0,0,0,0,15,65472,0,0,0,0,0,0,31,65408,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,127,65024,0,0,0,0,0,0,127,65024,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,1023,61440,0,0,0,0,0,0,1023,57344,0,0,0,0,0,0,2047,49152,0,0,0,
	0,0,0,4095,32768,0,0,0,0,0,0,8191,0,0,0,0,0,0,0,16383,0,0,0,0,0,0,0,32766,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,1,65520,0,0,0,0,0,0,3,65504,0,0,0,0,0,0,7,65472,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,15,65408,0,0,2032,0,0,0,31,65280,0,0,4080,0,0,0,63,65024,0,0,8160,0,0,0,127,64512,0,0,8160,0,0,0,255,63488,0,0,16352,0,0,0,255,61440,0,0,16320,0,
	0,0,511,57344,0,0,32704,0,0,0,1023,49152,0,0,32704,0,0,0,2047,49152,0,0,65408,0,0,0,4095,32768,0,0,65408,0,0,0,8191,0,0,1,65408,0,0,0,8190,0,0,3,65280,0,0,0,16380,0,0,7,65280,0,0,0,32760,0,0,7,65280,0,0,0,65520,0,0,15,65024,0,0,1,65520,0,0,31,65024,0,0,1,65504,0,0,127,65024,0,0,3,65472,0,0,1023,64512,0,0,7,65535,65535,65535,65535,64512,0,0,15,65535,65535,65535,65535,64512,0,0,31,65535,65535,65535,65535,63488,0,0,63,65535,65535,65535,65535,63488,0,
	0,63,65535,65535,65535,65535,63488,0,0,127,65535,65535,65535,65535,61440,0,0,255,65535,65535,65535,65535,61440,0,0,511,65535,65535,65535,65535,61440,0,0,1023,65535,65535,65535,65535,57344,0,0,1023,65535,65535,65535,65535,57344,0,0,2047,65535,65535,65535,65535,57344,0,0,4095,65535,65535,65535,65535,49152,0,0,4095,65535,65535,65535,65535,49152,0,0,4095,65535,65535,65535,65535,49152,0,0,4095,65535,65535,65535,65535,32768,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--3:3920:5199
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,4095,65520,0,0,0,0,0,0,16383,65534,0,0,0,0,0,0,65535,65535,0,0,0,0,0,3,65535,65535,49152,0,0,0,0,15,65535,65535,61440,0,0,0,0,31,65535,65535,63488,0,0,0,0,63,65535,65535,64512,0,0,0,0,255,65535,65535,64512,0,0,0,0,511,65535,65535,65024,0,0,0,0,1023,65471,65535,65280,0,0,0,0,1023,63488,65535,65408,0,0,0,0,2047,57344,16383,65408,0,0,
	0,0,4095,49152,4095,65472,0,0,0,0,8191,32768,1023,65504,0,0,0,0,8191,0,511,65504,0,0,0,0,16380,0,255,65520,0,0,0,0,32760,0,127,65520,0,0,0,0,32760,0,31,65528,0,0,0,0,65520,0,15,65528,0,0,0,1,65504,0,15,65532,0,0,0,1,65472,0,7,65532,0,0,0,1,65472,0,3,65532,0,0,0,3,65408,0,3,65532,0,0,0,3,65280,0,1,65534,0,0,0,7,65024,0,1,65534,0,0,0,7,65024,0,0,65534,0,0,0,15,64512,0,0,65534,0,0,0,15,64512,0,0,65534,0,0,
	0,15,63488,0,0,32766,0,0,0,31,61440,0,0,32766,0,0,0,31,61440,0,0,32766,0,0,0,31,57344,0,0,32766,0,0,0,31,57344,0,0,32766,0,0,0,63,49152,0,0,32766,0,0,0,63,32768,0,0,32766,0,0,0,63,32768,0,0,32766,0,0,0,1,0,0,0,32764,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,32760,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,0,65520,0,0,
	0,0,0,0,1,65520,0,0,0,0,0,0,1,65504,0,0,0,0,0,0,3,65504,0,0,0,0,0,0,7,65472,0,0,0,0,0,0,7,65408,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,127,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,1023,61440,0,0,0,0,0,0,2047,57344,0,0,0,0,0,0,4095,32768,0,0,0,0,0,0,8191,0,0,0,0,0,0,0,32766,0,0,0,
	0,0,0,0,65532,0,0,0,0,0,0,3,65534,0,0,0,0,0,0,7,65535,0,0,0,0,0,0,31,65535,49152,0,0,0,0,0,127,65535,61440,0,0,0,0,0,511,65535,63488,0,0,0,0,0,2047,65535,64512,0,0,0,0,0,8191,65535,65024,0,0,0,0,0,65535,65535,65280,0,0,0,0,3,65535,65535,65408,0,0,0,0,7,65535,65535,65472,0,0,0,0,7,65535,65535,65504,0,0,0,0,7,65535,65535,65520,0,0,0,0,7,65535,65535,65528,0,0,0,0,0,63,65535,65528,0,0,0,0,0,1,65535,65532,0,0,
	0,0,0,0,16383,65534,0,0,0,0,0,0,2047,65535,0,0,0,0,0,0,511,65535,32768,0,0,0,0,0,127,65535,32768,0,0,0,0,0,31,65535,49152,0,0,0,0,0,7,65535,49152,0,0,0,0,0,3,65535,57344,0,0,0,0,0,1,65535,57344,0,0,0,0,0,0,65535,61440,0,0,0,0,0,0,32767,61440,0,0,0,0,0,0,16383,61440,0,0,0,0,0,0,8191,61440,0,0,0,0,0,0,8191,63488,0,0,0,0,0,0,4095,63488,0,0,0,0,0,0,4095,63488,0,0,0,0,0,0,2047,63488,0,
	0,0,0,0,0,2047,63488,0,0,0,0,0,0,1023,64512,0,0,0,0,0,0,1023,64512,0,0,0,0,0,0,511,64512,0,0,0,0,0,0,511,64512,0,0,0,0,0,0,511,64512,0,0,0,0,0,0,511,64512,0,0,0,0,0,0,511,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,
	0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,61440,0,0,0,0,0,0,255,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,57344,0,0,0,0,0,0,511,57344,0,0,0,0,0,0,1023,49152,0,0,0,0,0,0,1023,49152,0,0,0,0,0,0,2047,49152,0,0,0,0,0,0,2047,32768,0,
	0,0,0,0,0,4095,32768,0,0,0,0,0,0,4095,0,0,0,0,0,0,0,8190,0,0,0,0,0,0,0,16382,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,32760,0,0,0,0,0,0,0,65520,0,0,0,0,0,0,3,65504,0,0,0,7,49152,0,7,65504,0,0,0,31,63488,0,15,65472,0,0,0,63,65024,0,31,65280,0,0,0,63,65408,0,127,65024,0,0,0,127,65520,0,255,64512,0,0,0,127,65532,0,2047,63488,0,0,0,127,65535,32768,8191,61440,0,0,0,127,65535,65031,65535,57344,0,0,
	0,127,65535,65535,65535,49152,0,0,0,127,65535,65535,65535,0,0,0,0,127,65535,65535,65534,0,0,0,0,127,65535,65535,65528,0,0,0,0,63,65535,65535,65520,0,0,0,0,63,65535,65535,65472,0,0,0,0,31,65535,65535,65280,0,0,0,0,7,65535,65535,64512,0,0,0,0,1,65535,65535,61440,0,0,0,0,0,32767,65535,32768,0,0,0,0,0,4095,65528,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--4:5200:6479
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,32512,0,0,0,0,0,0,0,65280,0,0,0,0,0,0,0,65280,0,0,0,0,0,0,1,65280,0,0,0,0,0,0,1,65280,0,0,0,0,0,0,3,65280,0,0,0,0,0,0,7,65280,0,0,0,0,0,0,7,65280,0,0,0,0,0,0,15,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,63,65280,0,0,
	0,0,0,0,63,65280,0,0,0,0,0,0,127,65280,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,511,65280,0,0,0,0,0,0,1023,65280,0,0,0,0,0,0,1023,65280,0,0,0,0,0,0,2047,65280,0,0,0,0,0,0,2047,65280,0,0,0,0,0,0,4095,65280,0,0,0,0,0,0,8191,65280,0,0,0,0,0,0,8191,65280,0,0,0,0,0,0,16383,65280,0,0,0,0,0,0,16383,65280,0,0,0,0,0,0,32767,65280,0,0,0,0,0,0,65535,65280,0,0,
	0,0,0,0,65471,65280,0,0,0,0,0,1,65471,65280,0,0,0,0,0,3,65343,65280,0,0,0,0,0,3,65343,65280,0,0,0,0,0,7,65087,65280,0,0,0,0,0,7,64575,65280,0,0,0,0,0,15,64575,65280,0,0,0,0,0,31,63551,65280,0,0,0,0,0,31,63551,65280,0,0,0,0,0,63,61503,65280,0,0,0,0,0,127,57407,65280,0,0,0,0,0,127,57407,65280,0,0,0,0,0,255,49215,65280,0,0,0,0,0,255,49215,65280,0,0,0,0,0,511,32831,65280,0,0,0,0,0,1023,63,65280,0,0,
	0,0,0,1023,63,65280,0,0,0,0,0,2046,63,65280,0,0,0,0,0,4094,63,65280,0,0,0,0,0,4092,63,65280,0,0,0,0,0,8184,63,65280,0,0,0,0,0,8184,63,65280,0,0,0,0,0,16368,63,65280,0,0,0,0,0,32752,63,65280,0,0,0,0,0,32736,63,65280,0,0,0,0,0,65472,63,65280,0,0,0,0,1,65472,63,65280,0,0,0,0,1,65408,63,65280,0,0,0,0,3,65408,63,65280,0,0,0,0,3,65280,63,65280,0,0,0,0,7,65024,63,65280,0,0,0,0,15,65024,63,65280,0,0,
	0,0,15,64512,63,65280,0,0,0,0,31,64512,63,65280,0,0,0,0,31,63488,63,65280,0,0,0,0,63,63488,63,65280,0,0,0,0,127,61440,63,65280,0,0,0,0,127,57344,63,65280,0,0,0,0,255,57344,63,65280,0,0,0,0,511,49152,63,65280,0,0,0,0,511,49152,63,65280,0,0,0,0,1023,32768,63,65280,0,0,0,0,1023,0,63,65280,0,0,0,0,2047,0,63,65280,0,0,0,0,4094,0,63,65280,0,0,0,0,4094,0,63,65280,0,0,0,0,8188,0,63,65280,0,0,0,0,16376,0,63,65280,0,0,
	0,0,16376,0,63,65280,0,0,0,0,32752,0,63,65280,0,0,0,0,32752,0,63,65280,0,0,0,0,65504,0,63,65280,0,0,0,1,65472,0,63,65280,0,0,0,1,65472,0,63,65280,0,0,0,3,65408,0,63,65280,0,0,0,7,65408,0,63,65280,0,0,0,7,65280,0,63,65280,0,0,0,15,65024,0,63,65280,0,0,0,15,65024,0,63,65280,0,0,0,31,64512,0,63,65280,0,0,0,63,64512,0,63,65280,0,0,0,63,63488,0,63,65280,0,0,0,127,63488,0,63,65280,0,0,0,255,61440,0,63,65280,0,0,
	0,255,57344,0,63,65280,0,0,0,511,57344,0,63,65280,0,0,0,511,49152,0,63,65280,0,0,0,1023,49152,0,63,65280,0,0,0,2047,32768,0,63,65280,0,0,0,2047,0,0,63,65280,0,0,0,4095,0,0,63,65280,0,0,0,8190,0,0,63,65280,0,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,
	0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,8191,65535,65535,65535,65535,65528,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,
	0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,
	0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--5:6480:7759
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,32512,0,0,0,0,0,0,0,65024,0,0,0,0,0,0,1,65024,0,0,0,0,0,0,7,65024,0,0,0,0,0,0,15,64512,0,0,0,0,0,0,127,64512,0,0,0,0,8191,65535,65535,64512,0,0,0,0,16383,65535,65535,63488,0,0,0,0,16383,65535,65535,63488,0,0,0,0,16383,65535,65535,63488,0,0,0,0,32767,65535,65535,61440,0,0,0,0,32767,65535,65535,61440,0,0,0,0,65535,65535,65535,57344,0,0,0,0,65535,65535,65535,57344,0,
	0,0,0,65535,65535,65535,57344,0,0,0,1,65535,65535,65535,49152,0,0,0,1,65535,65535,65535,49152,0,0,0,3,65535,65535,65535,49152,0,0,0,3,65535,65535,65535,32768,0,0,0,3,65535,65535,65535,32768,0,0,0,7,65535,65535,65534,0,0,0,0,7,65472,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,63,64512,0,0,0,0,
	0,0,127,64512,0,0,0,0,0,0,127,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,61440,0,0,0,0,0,0,255,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,57344,0,0,0,0,0,0,1023,57344,0,0,0,0,0,0,1023,49152,0,0,0,0,0,0,1023,49152,0,0,0,0,0,0,2047,32768,0,0,0,0,0,0,2047,32768,0,0,0,0,0,0,4095,0,0,0,0,0,0,0,4095,61440,0,0,0,0,0,0,4095,65024,0,0,0,0,0,0,8191,65504,0,0,0,0,
	0,0,8191,65532,0,0,0,0,0,0,16383,65535,32768,0,0,0,0,0,16383,65535,57344,0,0,0,0,0,16383,65535,63488,0,0,0,0,0,32767,65535,65024,0,0,0,0,0,32767,65535,65408,0,0,0,0,0,65535,65535,65504,0,0,0,0,0,65535,65535,65520,0,0,0,0,0,65535,65535,65532,0,0,0,0,1,65535,65535,65534,0,0,0,0,1,65535,65535,65535,0,0,0,0,3,65535,65535,65535,32768,0,0,0,3,65535,65535,65535,57344,0,0,0,3,65535,65535,65535,61440,0,0,0,3,65535,65535,65535,63488,0,0,0,3,65535,65535,65535,64512,0,0,
	0,0,32767,65535,65535,65024,0,0,0,0,15,65535,65535,65024,0,0,0,0,0,32767,65535,65280,0,0,0,0,0,2047,65535,65408,0,0,0,0,0,255,65535,65472,0,0,0,0,0,31,65535,65504,0,0,0,0,0,3,65535,65504,0,0,0,0,0,0,65535,65520,0,0,0,0,0,0,16383,65528,0,0,0,0,0,0,4095,65528,0,0,0,0,0,0,2047,65532,0,0,0,0,0,0,511,65534,0,0,0,0,0,0,255,65534,0,0,0,0,0,0,127,65534,0,0,0,0,0,0,31,65535,0,0,0,0,0,0,15,65535,0,0,
	0,0,0,0,7,65535,32768,0,0,0,0,0,3,65535,32768,0,0,0,0,0,3,65535,49152,0,0,0,0,0,1,65535,49152,0,0,0,0,0,0,65535,49152,0,0,0,0,0,0,32767,57344,0,0,0,0,0,0,32767,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,8191,57344,0,0,0,0,0,0,8191,61440,0,0,0,0,0,0,4095,61440,0,0,0,0,0,0,4095,61440,0,0,0,0,0,0,2047,61440,0,0,0,0,0,0,2047,61440,0,0,0,0,0,0,2047,63488,0,0,0,0,0,0,1023,63488,0,
	0,0,0,0,0,1023,63488,0,0,0,0,0,0,1023,63488,0,0,0,0,0,0,1023,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,511,63488,0,
	0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,57344,0,0,0,0,0,0,511,57344,0,0,0,0,0,0,511,57344,0,0,0,0,0,0,1023,57344,0,0,0,0,0,0,1023,49152,0,0,0,0,0,0,1023,49152,0,0,0,0,0,0,1023,32768,0,0,0,0,0,0,2047,32768,0,0,0,0,0,0,2047,32768,0,0,0,0,0,0,2047,0,0,0,0,0,0,0,4095,0,0,
	0,0,0,0,0,4094,0,0,0,0,0,0,0,4094,0,0,0,0,0,0,0,8188,0,0,0,0,0,0,0,8188,0,0,0,0,0,0,0,16376,0,0,0,0,0,0,0,16368,0,0,0,0,0,0,0,32752,0,0,0,0,0,0,0,65504,0,0,0,0,0,0,1,65472,0,0,0,0,0,0,1,65408,0,0,0,15,61440,0,3,65408,0,0,0,63,65280,0,15,65280,0,0,0,127,65504,0,31,65024,0,0,0,127,65528,0,63,64512,0,0,0,255,65535,0,255,63488,0,0,0,255,65535,49152,511,61440,0,0,
	0,255,65535,64512,4095,57344,0,0,0,255,65535,65472,32767,49152,0,0,0,255,65535,65535,65535,32768,0,0,0,255,65535,65535,65535,0,0,0,0,127,65535,65535,65534,0,0,0,0,127,65535,65535,65532,0,0,0,0,63,65535,65535,65520,0,0,0,0,31,65535,65535,65504,0,0,0,0,15,65535,65535,65408,0,0,0,0,7,65535,65535,65024,0,0,0,0,1,65535,65535,63488,0,0,0,0,0,65535,65535,49152,0,0,0,0,0,8191,65532,0,0,0,0,0,0,511,65408,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--6:7760:9039
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,64512,0,0,0,0,0,0,127,64512,0,0,0,0,0,0,4095,64512,0,0,0,0,0,0,32767,65024,0,0,0,0,0,3,65535,65024,0,0,0,0,0,31,65535,65024,0,0,0,0,0,127,65535,65024,0,0,0,0,0,511,65535,64512,0,0,0,0,0,2047,65535,49152,0,0,0,0,0,8191,65532,0,0,0,0,0,0,32767,65504,0,0,0,0,0,1,65535,65280,0,0,0,0,0,3,65535,64512,0,0,0,0,0,7,65535,57344,0,0,
	0,0,0,31,65535,32768,0,0,0,0,0,63,65534,0,0,0,0,0,0,127,65528,0,0,0,0,0,0,255,65520,0,0,0,0,0,0,511,65472,0,0,0,0,0,0,1023,65280,0,0,0,0,0,0,2047,65024,0,0,0,0,0,0,4095,64512,0,0,0,0,0,0,8191,61440,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,65535,32768,0,0,0,0,0,1,65534,0,0,0,0,0,0,1,65532,0,0,0,0,0,0,3,65528,0,0,0,0,0,0,7,65528,0,0,0,0,
	0,0,15,65520,0,0,0,0,0,0,31,65504,0,0,0,0,0,0,63,65472,0,0,0,0,0,0,127,65408,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,511,65024,0,0,0,0,0,0,1023,64512,0,0,0,0,0,0,2047,63488,0,0,0,0,0,0,2047,61440,0,0,0,0,0,0,4095,61440,0,0,0,0,0,0,8191,57344,0,0,0,0,0,0,8191,57344,0,0,0,0,0,0,16383,49152,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,32767,32768,0,0,0,0,
	0,0,65535,0,0,0,0,0,0,1,65535,0,0,0,0,0,0,1,65534,0,0,0,0,0,0,3,65534,0,0,0,0,0,0,3,65534,0,0,0,0,0,0,3,65532,0,0,0,0,0,0,7,65532,0,0,0,0,0,0,7,65528,0,0,0,0,0,0,15,65528,0,0,0,0,0,0,15,65528,7,65532,0,0,0,0,31,65520,127,65535,32768,0,0,0,31,65520,511,65535,61440,0,0,0,63,65520,4095,65535,64512,0,0,0,63,65504,8191,65535,65024,0,0,0,63,65504,32767,65535,65408,0,0,0,127,65504,65535,65535,65472,0,0,
	0,127,65507,65535,65535,65504,0,0,0,127,65511,65535,65535,65520,0,0,0,255,65487,65535,65535,65528,0,0,0,255,65503,65535,65535,65532,0,0,0,255,65503,65535,65535,65534,0,0,0,255,65535,65532,8191,65535,0,0,0,511,65535,65024,255,65535,32768,0,0,511,65535,61440,63,65535,49152,0,0,511,65535,49152,15,65535,49152,0,0,511,65535,0,7,65535,57344,0,0,511,65532,0,1,65535,61440,0,0,1023,65528,0,0,65535,61440,0,0,1023,65520,0,0,32767,63488,0,0,1023,65504,0,0,32767,63488,0,0,1023,65408,0,0,16383,64512,0,0,1023,65408,0,0,8191,64512,0,
	0,1023,65280,0,0,4095,65024,0,0,1023,65280,0,0,4095,65024,0,0,1023,65024,0,0,2047,65024,0,0,1023,65024,0,0,2047,65280,0,0,2047,65024,0,0,1023,65280,0,0,2047,64512,0,0,1023,65280,0,0,2047,64512,0,0,1023,65408,0,0,2047,64512,0,0,511,65408,0,0,2047,64512,0,0,511,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65472,0,0,2047,63488,0,0,255,65472,0,0,2047,63488,0,0,127,65472,0,0,2047,63488,0,0,127,65472,0,0,2047,63488,0,0,127,65472,0,
	0,2047,63488,0,0,127,65472,0,0,2047,63488,0,0,63,65504,0,0,1023,63488,0,0,63,65504,0,0,1023,63488,0,0,63,65504,0,0,1023,63488,0,0,63,65504,0,0,1023,63488,0,0,63,65504,0,0,1023,63488,0,0,63,65504,0,0,1023,63488,0,0,63,65504,0,0,1023,64512,0,0,31,65504,0,0,1023,64512,0,0,31,65504,0,0,1023,64512,0,0,31,65504,0,0,1023,64512,0,0,31,65504,0,0,511,64512,0,0,31,65504,0,0,511,64512,0,0,31,65504,0,0,511,64512,0,0,31,65504,0,0,511,64512,0,0,31,65504,0,
	0,511,64512,0,0,31,65504,0,0,511,65024,0,0,31,65504,0,0,255,65024,0,0,31,65472,0,0,255,65024,0,0,31,65472,0,0,255,65024,0,0,31,65472,0,0,255,65024,0,0,31,65472,0,0,255,65024,0,0,31,65472,0,0,127,65280,0,0,31,65472,0,0,127,65280,0,0,31,65408,0,0,127,65280,0,0,31,65408,0,0,63,65408,0,0,63,65408,0,0,63,65408,0,0,63,65408,0,0,63,65408,0,0,63,65280,0,0,63,65472,0,0,63,65280,0,0,31,65472,0,0,63,65280,0,0,31,65472,0,0,127,65024,0,
	0,15,65504,0,0,127,65024,0,0,15,65504,0,0,127,65024,0,0,15,65520,0,0,127,64512,0,0,7,65520,0,0,255,64512,0,0,7,65528,0,0,255,63488,0,0,3,65528,0,0,255,63488,0,0,3,65532,0,0,511,61440,0,0,1,65532,0,0,511,61440,0,0,1,65534,0,0,1023,61440,0,0,0,65534,0,0,2047,57344,0,0,0,32767,0,0,2047,49152,0,0,0,32767,32768,0,4095,49152,0,0,0,16383,57344,0,8191,32768,0,0,0,8191,61440,0,32767,0,0,0,0,8191,63488,0,65535,0,0,0,0,4095,65024,1,65534,0,0,
	0,0,2047,65280,7,65532,0,0,0,0,1023,65504,63,65528,0,0,0,0,511,65535,1023,65520,0,0,0,0,255,65535,65535,65504,0,0,0,0,127,65535,65535,65472,0,0,0,0,63,65535,65535,65408,0,0,0,0,15,65535,65535,65024,0,0,0,0,7,65535,65535,64512,0,0,0,0,1,65535,65535,61440,0,0,0,0,0,32767,65535,49152,0,0,0,0,0,8191,65535,0,0,0,0,0,0,1023,65528,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--7:9040:10319
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,65535,65535,65535,65535,65472,0,0,0,65535,65535,65535,65535,65472,0,0,1,65535,65535,65535,65535,65472,0,0,1,65535,65535,65535,65535,65472,0,0,1,65535,65535,65535,65535,65472,0,0,1,65535,65535,65535,65535,65408,0,0,3,65535,65535,65535,65535,65408,0,0,3,65535,65535,65535,65535,65408,0,0,3,65535,65535,65535,65535,65408,0,0,7,65535,65535,65535,65535,65280,0,0,7,65535,65535,65535,65535,65280,0,
	0,7,65535,65535,65535,65535,65280,0,0,15,65535,65535,65535,65535,65024,0,0,15,65535,65535,65535,65535,65024,0,0,15,65528,0,0,31,65024,0,0,31,65472,0,0,31,65024,0,0,31,65280,0,0,63,64512,0,0,31,65024,0,0,63,64512,0,0,63,64512,0,0,63,64512,0,0,63,63488,0,0,63,63488,0,0,63,63488,0,0,127,63488,0,0,127,61440,0,0,127,63488,0,0,127,61440,0,0,127,63488,0,0,127,57344,0,0,255,61440,0,0,255,49152,0,0,255,61440,0,0,255,49152,0,0,255,61440,0,0,255,32768,0,0,511,57344,0,
	0,511,32768,0,0,511,57344,0,0,511,0,0,0,511,57344,0,0,1023,0,0,0,511,57344,0,0,1022,0,0,0,1023,49152,0,0,1020,0,0,0,1023,49152,0,0,2044,0,0,0,1023,49152,0,0,1016,0,0,0,2047,32768,0,0,0,0,0,0,2047,32768,0,0,0,0,0,0,2047,32768,0,0,0,0,0,0,4095,32768,0,0,0,0,0,0,4095,0,0,0,0,0,0,0,4095,0,0,0,0,0,0,0,8191,0,0,0,0,0,0,0,8191,0,0,0,0,0,0,0,8190,0,0,0,0,0,0,0,8190,0,0,
	0,0,0,0,0,16382,0,0,0,0,0,0,0,16380,0,0,0,0,0,0,0,16380,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,32760,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,0,65520,0,0,0,0,0,0,0,65520,0,0,0,0,0,0,1,65520,0,0,0,0,0,0,1,65520,0,0,0,0,0,0,1,65504,0,0,0,0,0,0,3,65504,0,0,0,0,0,0,3,65504,0,0,0,0,0,0,3,65472,0,0,
	0,0,0,0,7,65472,0,0,0,0,0,0,7,65472,0,0,0,0,0,0,7,65472,0,0,0,0,0,0,7,65408,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,15,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,31,65280,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,63,64512,0,0,0,0,0,0,127,64512,0,0,0,0,0,0,127,64512,0,0,
	0,0,0,0,127,64512,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,255,63488,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,511,61440,0,0,0,0,0,0,1023,57344,0,0,0,0,0,0,1023,57344,0,0,0,0,0,0,1023,57344,0,0,0,0,0,0,2047,49152,0,0,0,0,0,0,2047,49152,0,0,0,0,0,0,2047,49152,0,0,0,0,0,0,4095,49152,0,0,0,0,0,0,4095,32768,0,0,
	0,0,0,0,4095,32768,0,0,0,0,0,0,8191,32768,0,0,0,0,0,0,8191,32768,0,0,0,0,0,0,8191,0,0,0,0,0,0,0,8191,0,0,0,0,0,0,0,16383,0,0,0,0,0,0,0,16382,0,0,0,0,0,0,0,16382,0,0,0,0,0,0,0,32766,0,0,0,0,0,0,0,32766,0,0,0,0,0,0,0,32764,0,0,0,0,0,0,0,65532,0,0,0,0,0,0,0,65532,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,0,65528,0,0,0,0,0,0,1,65528,0,0,0,
	0,0,0,1,65528,0,0,0,0,0,0,1,65520,0,0,0,0,0,0,3,65520,0,0,0,0,0,0,3,65520,0,0,0,0,0,0,3,65504,0,0,0,0,0,0,7,65504,0,0,0,0,0,0,7,65504,0,0,0,0,0,0,7,65504,0,0,0,0,0,0,7,65472,0,0,0,0,0,0,15,65472,0,0,0,0,0,0,15,65472,0,0,0,0,0,0,15,65408,0,0,0,0,0,0,31,65408,0,0,0,0,0,0,31,65408,0,0,0,0,0,0,31,65408,0,0,0,0,0,0,63,65280,0,0,0,
	0,0,0,63,65280,0,0,0,0,0,0,63,65280,0,0,0,0,0,0,63,65024,0,0,0,0,0,0,127,65024,0,0,0,0,0,0,127,65024,0,0,0,0,0,0,127,65024,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,255,64512,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,511,63488,0,0,0,0,0,0,1023,63488,0,0,0,0,0,0,1023,61440,0,0,0,0,0,0,1023,61440,0,0,0,0,0,0,1023,61440,0,0,0,
	0,0,0,2047,57344,0,0,0,0,0,0,2047,57344,0,0,0,0,0,0,2047,57344,0,0,0,0,0,0,4095,57344,0,0,0,0,0,0,4095,49152,0,0,0,0,0,0,4095,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,8191,49152,0,0,0,0,0,0,8191,32768,0,0,0,0,0,0,8191,32768,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--8:10320:11599
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,255,65280,0,0,0,0,0,0,4095,65520,0,0,0,0,0,0,32767,65534,0,0,0,0,0,1,65535,65535,32768,0,0,0,0,7,65535,65535,57344,0,0,0,0,31,65535,65535,63488,0,0,0,0,63,65535,65535,64512,0,0,0,0,255,65535,65535,65024,0,0,0,0,511,65535,65535,65408,0,0,0,0,1023,65520,65535,65472,0,0,0,0,2047,64512,1023,65504,0,0,0,0,4095,57344,127,65504,0,0,0,0,8191,32768,15,65520,0,0,
	0,0,16383,0,7,65528,0,0,0,0,32764,0,1,65532,0,0,0,0,65528,0,0,65532,0,0,0,0,65520,0,0,32766,0,0,0,1,65520,0,0,32766,0,0,0,3,65504,0,0,16383,0,0,0,3,65472,0,0,8191,0,0,0,7,65408,0,0,8191,32768,0,0,7,65408,0,0,4095,32768,0,0,7,65408,0,0,4095,32768,0,0,15,65280,0,0,4095,49152,0,0,15,65280,0,0,2047,49152,0,0,15,65280,0,0,2047,49152,0,0,31,65024,0,0,2047,49152,0,0,31,65024,0,0,2047,49152,0,0,31,65024,0,0,2047,49152,0,
	0,31,65024,0,0,2047,49152,0,0,31,65024,0,0,2047,57344,0,0,31,65280,0,0,2047,57344,0,0,31,65280,0,0,2047,57344,0,0,63,65280,0,0,2047,49152,0,0,63,65280,0,0,2047,49152,0,0,63,65280,0,0,2047,49152,0,0,63,65280,0,0,2047,49152,0,0,31,65408,0,0,2047,49152,0,0,31,65408,0,0,4095,49152,0,0,31,65408,0,0,4095,49152,0,0,31,65472,0,0,4095,32768,0,0,31,65472,0,0,4095,32768,0,0,31,65504,0,0,8191,32768,0,0,31,65504,0,0,8191,32768,0,0,31,65520,0,0,8191,0,0,
	0,15,65528,0,0,16383,0,0,0,15,65528,0,0,16382,0,0,0,15,65532,0,0,32766,0,0,0,15,65534,0,0,32764,0,0,0,7,65535,0,0,65532,0,0,0,7,65535,32768,1,65532,0,0,0,7,65535,32768,1,65528,0,0,0,3,65535,49152,3,65520,0,0,0,3,65535,57344,7,65504,0,0,0,1,65535,61440,15,65504,0,0,0,0,65535,64512,31,65472,0,0,0,0,65535,65024,63,65408,0,0,0,0,32767,65280,127,65280,0,0,0,0,16383,65408,255,65024,0,0,0,0,16383,65504,511,64512,0,0,0,0,8191,65520,1023,63488,0,0,
	0,0,4095,65532,2047,61440,0,0,0,0,2047,65534,8191,57344,0,0,0,0,1023,65535,49151,32768,0,0,0,0,511,65535,65535,0,0,0,0,0,255,65535,65532,0,0,0,0,0,127,65535,65528,0,0,0,0,0,63,65535,65504,0,0,0,0,0,31,65535,65408,0,0,0,0,0,15,65535,65408,0,0,0,0,0,7,65535,65472,0,0,0,0,0,3,65535,65504,0,0,0,0,0,1,65535,65528,0,0,0,0,0,0,65535,65532,0,0,0,0,0,0,32767,65534,0,0,0,0,0,0,16383,65535,32768,0,0,0,0,0,16383,65535,49152,0,0,
	0,0,0,65535,65535,57344,0,0,0,0,1,65535,65535,61440,0,0,0,0,3,65535,65535,63488,0,0,0,0,7,65535,65535,64512,0,0,0,0,31,65487,65535,65024,0,0,0,0,63,65415,65535,65280,0,0,0,0,127,65283,65535,65408,0,0,0,0,255,65024,65535,65472,0,0,0,0,511,64512,32767,65504,0,0,0,0,1023,63488,8191,65520,0,0,0,0,2047,61440,4095,65528,0,0,0,0,4095,57344,2047,65532,0,0,0,0,8191,49152,1023,65532,0,0,0,0,16383,32768,255,65534,0,0,0,0,32767,0,127,65534,0,0,0,0,32766,0,63,65535,0,0,
	0,0,65532,0,31,65535,32768,0,0,1,65528,0,15,65535,32768,0,0,1,65528,0,7,65535,49152,0,0,3,65520,0,3,65535,49152,0,0,3,65520,0,1,65535,57344,0,0,7,65504,0,0,65535,57344,0,0,7,65504,0,0,32767,61440,0,0,15,65472,0,0,16383,61440,0,0,15,65472,0,0,8191,61440,0,0,15,65408,0,0,8191,63488,0,0,31,65408,0,0,4095,63488,0,0,31,65408,0,0,2047,63488,0,0,31,65280,0,0,2047,63488,0,0,31,65280,0,0,1023,64512,0,0,63,65280,0,0,1023,64512,0,0,63,65280,0,0,511,64512,0,
	0,63,65280,0,0,511,64512,0,0,63,65024,0,0,511,64512,0,0,63,65024,0,0,255,64512,0,0,63,65024,0,0,255,64512,0,0,63,65024,0,0,255,64512,0,0,63,65024,0,0,255,64512,0,0,127,65024,0,0,127,64512,0,0,127,65024,0,0,127,64512,0,0,127,65024,0,0,127,64512,0,0,127,65024,0,0,127,64512,0,0,63,65280,0,0,127,64512,0,0,63,65280,0,0,127,64512,0,0,63,65280,0,0,127,64512,0,0,63,65280,0,0,127,64512,0,0,63,65280,0,0,127,64512,0,0,63,65280,0,0,127,64512,0,
	0,31,65408,0,0,127,63488,0,0,31,65408,0,0,127,63488,0,0,31,65408,0,0,127,63488,0,0,15,65472,0,0,255,63488,0,0,15,65472,0,0,255,61440,0,0,15,65472,0,0,255,61440,0,0,7,65504,0,0,511,57344,0,0,7,65520,0,0,511,57344,0,0,3,65520,0,0,1023,49152,0,0,1,65528,0,0,1023,49152,0,0,1,65532,0,0,2047,32768,0,0,0,65534,0,0,4095,32768,0,0,0,32767,0,0,8191,0,0,0,0,32767,32768,0,16382,0,0,0,0,16383,57344,0,65534,0,0,0,0,8191,63488,1,65532,0,0,
	0,0,4095,65024,15,65528,0,0,0,0,2047,65472,127,65520,0,0,0,0,1023,65535,49151,65504,0,0,0,0,511,65535,65535,65472,0,0,0,0,255,65535,65535,65408,0,0,0,0,127,65535,65535,65024,0,0,0,0,31,65535,65535,64512,0,0,0,0,15,65535,65535,61440,0,0,0,0,3,65535,65535,49152,0,0,0,0,0,65535,65534,0,0,0,0,0,0,4095,65520,0,0,0,0,0,0,255,65024,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--9:11600:12879
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1023,64512,0,0,0,0,0,0,16383,65472,0,0,0,0,0,0,65535,65520,0,0,0,0,0,3,65535,65532,0,0,0,0,0,15,65535,65535,0,0,0,0,0,63,65535,65535,49152,0,0,0,0,127,65535,65535,57344,0,0,0,0,255,65535,65535,61440,0,0,0,0,1023,65408,32767,64512,0,0,0,0,2047,64512,4095,65024,0,0,0,0,4095,61440,1023,65280,0,0,0,0,8191,49152,255,65408,0,0,0,0,8191,32768,127,65472,0,0,0,0,16383,0,63,65504,0,0,
	0,0,32766,0,31,65504,0,0,0,0,65532,0,15,65520,0,0,0,0,65532,0,7,65528,0,0,0,1,65528,0,3,65532,0,0,0,1,65520,0,3,65532,0,0,0,3,65504,0,1,65534,0,0,0,7,65504,0,0,65534,0,0,0,7,65472,0,0,65535,0,0,0,15,65472,0,0,32767,32768,0,0,31,65408,0,0,32767,32768,0,0,31,65408,0,0,16383,49152,0,0,31,65408,0,0,16383,49152,0,0,63,65280,0,0,16383,57344,0,0,63,65280,0,0,8191,57344,0,0,63,65280,0,0,8191,61440,0,0,127,65024,0,0,4095,61440,0,
	0,127,65024,0,0,4095,61440,0,0,255,65024,0,0,4095,63488,0,0,255,65024,0,0,4095,63488,0,0,255,64512,0,0,2047,63488,0,0,255,64512,0,0,2047,64512,0,0,511,64512,0,0,2047,64512,0,0,511,64512,0,0,1023,64512,0,0,511,64512,0,0,1023,65024,0,0,511,64512,0,0,1023,65024,0,0,1023,64512,0,0,1023,65024,0,0,1023,64512,0,0,1023,65024,0,0,1023,63488,0,0,511,65024,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,
	0,1023,63488,0,0,255,65280,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,127,65408,0,0,2047,64512,0,0,127,65408,0,0,1023,65024,0,0,127,65472,0,0,1023,65024,0,0,127,65472,0,0,1023,65024,0,0,127,65472,0,
	0,1023,65024,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,511,65280,0,0,127,65472,0,0,511,65408,0,0,127,65408,0,0,511,65408,0,0,127,65408,0,0,511,65472,0,0,127,65408,0,0,255,65472,0,0,127,65408,0,0,255,65472,0,0,127,65408,0,0,255,65504,0,0,127,65408,0,0,127,65504,0,0,127,65408,0,0,127,65520,0,0,255,65408,0,0,127,65528,0,0,255,65408,0,0,63,65528,0,0,255,65408,0,0,63,65532,0,0,511,65408,0,
	0,31,65534,0,0,1023,65408,0,0,31,65534,0,0,2047,65280,0,0,15,65535,0,0,4095,65280,0,0,15,65535,32768,0,8191,65280,0,0,7,65535,57344,0,32767,65280,0,0,3,65535,61440,1,65535,65280,0,0,3,65535,64512,7,65535,65280,0,0,1,65535,65280,31,65535,65024,0,0,0,65535,65472,255,65535,65024,0,0,0,32767,65534,2047,65535,65024,0,0,0,16383,65535,65535,65023,65024,0,0,0,8191,65535,65535,63999,64512,0,0,0,4095,65535,65535,58367,64512,0,0,0,2047,65535,65535,50175,64512,0,0,0,511,65535,65535,1023,64512,0,0,0,255,65535,65532,2047,63488,0,
	0,0,63,65535,65520,2047,63488,0,0,0,15,65535,65280,2047,63488,0,0,0,1,65535,61440,4095,61440,0,0,0,0,992,0,4095,61440,0,0,0,0,0,0,8191,61440,0,0,0,0,0,0,8191,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,65535,32768,0,0,0,0,0,0,65535,32768,0,0,0,0,0,1,65535,0,0,0,0,0,0,3,65535,0,0,0,0,0,0,3,65534,0,0,0,0,0,0,7,65534,0,0,
	0,0,0,0,7,65534,0,0,0,0,0,0,15,65532,0,0,0,0,0,0,31,65528,0,0,0,0,0,0,31,65528,0,0,0,0,0,0,63,65520,0,0,0,0,0,0,127,65520,0,0,0,0,0,0,127,65504,0,0,0,0,0,0,255,65472,0,0,0,0,0,0,511,65472,0,0,0,0,0,0,1023,65408,0,0,0,0,0,0,1023,65280,0,0,0,0,0,0,2047,65280,0,0,0,0,0,0,4095,65024,0,0,0,0,0,0,8191,64512,0,0,0,0,0,0,16383,64512,0,0,0,0,0,0,32767,63488,0,0,
	0,0,0,0,32767,61440,0,0,0,0,0,0,65535,57344,0,0,0,0,0,3,65535,49152,0,0,0,0,0,7,65535,32768,0,0,0,0,0,15,65535,0,0,0,0,0,0,31,65534,0,0,0,0,0,0,63,65532,0,0,0,0,0,0,127,65528,0,0,0,0,0,0,511,65520,0,0,0,0,0,0,1023,65504,0,0,0,0,0,0,2047,65472,0,0,0,0,0,0,8191,65408,0,0,0,0,0,0,16383,65024,0,0,0,0,0,0,65535,64512,0,0,0,0,0,3,65535,63488,0,0,0,0,0,15,65535,57344,0,0,0,
	0,0,63,65535,49152,0,0,0,0,0,255,65535,0,0,0,0,0,0,1023,65532,0,0,0,0,0,0,8191,65528,0,0,0,0,0,0,65535,65504,0,0,0,0,0,15,65535,65408,0,0,0,0,0,63,65535,64512,0,0,0,0,0,63,65535,61440,0,0,0,0,0,63,65535,32768,0,0,0,0,0,63,65532,0,0,0,0,0,0,31,65472,0,0,0,0,0,0,31,63488,0,0,0,0,0,0,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--xx:補齊944空位
	--12880~16384-12880=3504-1280x2=944
	--1280
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1023,64512,0,0,0,0,0,0,16383,65472,0,0,0,0,0,0,65535,65520,0,0,0,0,0,3,65535,65532,0,0,0,0,0,15,65535,65535,0,0,0,0,0,63,65535,65535,49152,0,0,0,0,127,65535,65535,57344,0,0,0,0,255,65535,65535,61440,0,0,0,0,1023,65408,32767,64512,0,0,0,0,2047,64512,4095,65024,0,0,0,0,4095,61440,1023,65280,0,0,0,0,8191,49152,255,65408,0,0,0,0,8191,32768,127,65472,0,0,0,0,16383,0,63,65504,0,0,
	0,0,32766,0,31,65504,0,0,0,0,65532,0,15,65520,0,0,0,0,65532,0,7,65528,0,0,0,1,65528,0,3,65532,0,0,0,1,65520,0,3,65532,0,0,0,3,65504,0,1,65534,0,0,0,7,65504,0,0,65534,0,0,0,7,65472,0,0,65535,0,0,0,15,65472,0,0,32767,32768,0,0,31,65408,0,0,32767,32768,0,0,31,65408,0,0,16383,49152,0,0,31,65408,0,0,16383,49152,0,0,63,65280,0,0,16383,57344,0,0,63,65280,0,0,8191,57344,0,0,63,65280,0,0,8191,61440,0,0,127,65024,0,0,4095,61440,0,
	0,127,65024,0,0,4095,61440,0,0,255,65024,0,0,4095,63488,0,0,255,65024,0,0,4095,63488,0,0,255,64512,0,0,2047,63488,0,0,255,64512,0,0,2047,64512,0,0,511,64512,0,0,2047,64512,0,0,511,64512,0,0,1023,64512,0,0,511,64512,0,0,1023,65024,0,0,511,64512,0,0,1023,65024,0,0,1023,64512,0,0,1023,65024,0,0,1023,64512,0,0,1023,65024,0,0,1023,63488,0,0,511,65024,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,
	0,1023,63488,0,0,255,65280,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,127,65408,0,0,2047,64512,0,0,127,65408,0,0,1023,65024,0,0,127,65472,0,0,1023,65024,0,0,127,65472,0,0,1023,65024,0,0,127,65472,0,
	0,1023,65024,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,511,65280,0,0,127,65472,0,0,511,65408,0,0,127,65408,0,0,511,65408,0,0,127,65408,0,0,511,65472,0,0,127,65408,0,0,255,65472,0,0,127,65408,0,0,255,65472,0,0,127,65408,0,0,255,65504,0,0,127,65408,0,0,127,65504,0,0,127,65408,0,0,127,65520,0,0,255,65408,0,0,127,65528,0,0,255,65408,0,0,63,65528,0,0,255,65408,0,0,63,65532,0,0,511,65408,0,
	0,31,65534,0,0,1023,65408,0,0,31,65534,0,0,2047,65280,0,0,15,65535,0,0,4095,65280,0,0,15,65535,32768,0,8191,65280,0,0,7,65535,57344,0,32767,65280,0,0,3,65535,61440,1,65535,65280,0,0,3,65535,64512,7,65535,65280,0,0,1,65535,65280,31,65535,65024,0,0,0,65535,65472,255,65535,65024,0,0,0,32767,65534,2047,65535,65024,0,0,0,16383,65535,65535,65023,65024,0,0,0,8191,65535,65535,63999,64512,0,0,0,4095,65535,65535,58367,64512,0,0,0,2047,65535,65535,50175,64512,0,0,0,511,65535,65535,1023,64512,0,0,0,255,65535,65532,2047,63488,0,
	0,0,63,65535,65520,2047,63488,0,0,0,15,65535,65280,2047,63488,0,0,0,1,65535,61440,4095,61440,0,0,0,0,992,0,4095,61440,0,0,0,0,0,0,8191,61440,0,0,0,0,0,0,8191,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,65535,32768,0,0,0,0,0,0,65535,32768,0,0,0,0,0,1,65535,0,0,0,0,0,0,3,65535,0,0,0,0,0,0,3,65534,0,0,0,0,0,0,7,65534,0,0,
	0,0,0,0,7,65534,0,0,0,0,0,0,15,65532,0,0,0,0,0,0,31,65528,0,0,0,0,0,0,31,65528,0,0,0,0,0,0,63,65520,0,0,0,0,0,0,127,65520,0,0,0,0,0,0,127,65504,0,0,0,0,0,0,255,65472,0,0,0,0,0,0,511,65472,0,0,0,0,0,0,1023,65408,0,0,0,0,0,0,1023,65280,0,0,0,0,0,0,2047,65280,0,0,0,0,0,0,4095,65024,0,0,0,0,0,0,8191,64512,0,0,0,0,0,0,16383,64512,0,0,0,0,0,0,32767,63488,0,0,
	0,0,0,0,32767,61440,0,0,0,0,0,0,65535,57344,0,0,0,0,0,3,65535,49152,0,0,0,0,0,7,65535,32768,0,0,0,0,0,15,65535,0,0,0,0,0,0,31,65534,0,0,0,0,0,0,63,65532,0,0,0,0,0,0,127,65528,0,0,0,0,0,0,511,65520,0,0,0,0,0,0,1023,65504,0,0,0,0,0,0,2047,65472,0,0,0,0,0,0,8191,65408,0,0,0,0,0,0,16383,65024,0,0,0,0,0,0,65535,64512,0,0,0,0,0,3,65535,63488,0,0,0,0,0,15,65535,57344,0,0,0,
	0,0,63,65535,49152,0,0,0,0,0,255,65535,0,0,0,0,0,0,1023,65532,0,0,0,0,0,0,8191,65528,0,0,0,0,0,0,65535,65504,0,0,0,0,0,15,65535,65408,0,0,0,0,0,63,65535,64512,0,0,0,0,0,63,65535,61440,0,0,0,0,0,63,65535,32768,0,0,0,0,0,63,65532,0,0,0,0,0,0,31,65472,0,0,0,0,0,0,31,63488,0,0,0,0,0,0,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	--1280
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1023,64512,0,0,0,0,0,0,16383,65472,0,0,0,0,0,0,65535,65520,0,0,0,0,0,3,65535,65532,0,0,0,0,0,15,65535,65535,0,0,0,0,0,63,65535,65535,49152,0,0,0,0,127,65535,65535,57344,0,0,0,0,255,65535,65535,61440,0,0,0,0,1023,65408,32767,64512,0,0,0,0,2047,64512,4095,65024,0,0,0,0,4095,61440,1023,65280,0,0,0,0,8191,49152,255,65408,0,0,0,0,8191,32768,127,65472,0,0,0,0,16383,0,63,65504,0,0,
	0,0,32766,0,31,65504,0,0,0,0,65532,0,15,65520,0,0,0,0,65532,0,7,65528,0,0,0,1,65528,0,3,65532,0,0,0,1,65520,0,3,65532,0,0,0,3,65504,0,1,65534,0,0,0,7,65504,0,0,65534,0,0,0,7,65472,0,0,65535,0,0,0,15,65472,0,0,32767,32768,0,0,31,65408,0,0,32767,32768,0,0,31,65408,0,0,16383,49152,0,0,31,65408,0,0,16383,49152,0,0,63,65280,0,0,16383,57344,0,0,63,65280,0,0,8191,57344,0,0,63,65280,0,0,8191,61440,0,0,127,65024,0,0,4095,61440,0,
	0,127,65024,0,0,4095,61440,0,0,255,65024,0,0,4095,63488,0,0,255,65024,0,0,4095,63488,0,0,255,64512,0,0,2047,63488,0,0,255,64512,0,0,2047,64512,0,0,511,64512,0,0,2047,64512,0,0,511,64512,0,0,1023,64512,0,0,511,64512,0,0,1023,65024,0,0,511,64512,0,0,1023,65024,0,0,1023,64512,0,0,1023,65024,0,0,1023,64512,0,0,1023,65024,0,0,1023,63488,0,0,511,65024,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,0,1023,63488,0,0,511,65280,0,
	0,1023,63488,0,0,255,65280,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,63488,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,255,65408,0,0,2047,64512,0,0,127,65408,0,0,2047,64512,0,0,127,65408,0,0,1023,65024,0,0,127,65472,0,0,1023,65024,0,0,127,65472,0,0,1023,65024,0,0,127,65472,0,
	0,1023,65024,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,1023,65280,0,0,127,65472,0,0,511,65280,0,0,127,65472,0,0,511,65408,0,0,127,65408,0,0,511,65408,0,0,127,65408,0,0,511,65472,0,0,127,65408,0,0,255,65472,0,0,127,65408,0,0,255,65472,0,0,127,65408,0,0,255,65504,0,0,127,65408,0,0,127,65504,0,0,127,65408,0,0,127,65520,0,0,255,65408,0,0,127,65528,0,0,255,65408,0,0,63,65528,0,0,255,65408,0,0,63,65532,0,0,511,65408,0,
	0,31,65534,0,0,1023,65408,0,0,31,65534,0,0,2047,65280,0,0,15,65535,0,0,4095,65280,0,0,15,65535,32768,0,8191,65280,0,0,7,65535,57344,0,32767,65280,0,0,3,65535,61440,1,65535,65280,0,0,3,65535,64512,7,65535,65280,0,0,1,65535,65280,31,65535,65024,0,0,0,65535,65472,255,65535,65024,0,0,0,32767,65534,2047,65535,65024,0,0,0,16383,65535,65535,65023,65024,0,0,0,8191,65535,65535,63999,64512,0,0,0,4095,65535,65535,58367,64512,0,0,0,2047,65535,65535,50175,64512,0,0,0,511,65535,65535,1023,64512,0,0,0,255,65535,65532,2047,63488,0,
	0,0,63,65535,65520,2047,63488,0,0,0,15,65535,65280,2047,63488,0,0,0,1,65535,61440,4095,61440,0,0,0,0,992,0,4095,61440,0,0,0,0,0,0,8191,61440,0,0,0,0,0,0,8191,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,16383,57344,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,32767,49152,0,0,0,0,0,0,65535,32768,0,0,0,0,0,0,65535,32768,0,0,0,0,0,1,65535,0,0,0,0,0,0,3,65535,0,0,0,0,0,0,3,65534,0,0,0,0,0,0,7,65534,0,0,
	0,0,0,0,7,65534,0,0,0,0,0,0,15,65532,0,0,0,0,0,0,31,65528,0,0,0,0,0,0,31,65528,0,0,0,0,0,0,63,65520,0,0,0,0,0,0,127,65520,0,0,0,0,0,0,127,65504,0,0,0,0,0,0,255,65472,0,0,0,0,0,0,511,65472,0,0,0,0,0,0,1023,65408,0,0,0,0,0,0,1023,65280,0,0,0,0,0,0,2047,65280,0,0,0,0,0,0,4095,65024,0,0,0,0,0,0,8191,64512,0,0,0,0,0,0,16383,64512,0,0,0,0,0,0,32767,63488,0,0,
	0,0,0,0,32767,61440,0,0,0,0,0,0,65535,57344,0,0,0,0,0,3,65535,49152,0,0,0,0,0,7,65535,32768,0,0,0,0,0,15,65535,0,0,0,0,0,0,31,65534,0,0,0,0,0,0,63,65532,0,0,0,0,0,0,127,65528,0,0,0,0,0,0,511,65520,0,0,0,0,0,0,1023,65504,0,0,0,0,0,0,2047,65472,0,0,0,0,0,0,8191,65408,0,0,0,0,0,0,16383,65024,0,0,0,0,0,0,65535,64512,0,0,0,0,0,3,65535,63488,0,0,0,0,0,15,65535,57344,0,0,0,
	0,0,63,65535,49152,0,0,0,0,0,255,65535,0,0,0,0,0,0,1023,65532,0,0,0,0,0,0,8191,65528,0,0,0,0,0,0,65535,65504,0,0,0,0,0,15,65535,65408,0,0,0,0,0,63,65535,64512,0,0,0,0,0,63,65535,61440,0,0,0,0,0,63,65535,32768,0,0,0,0,0,63,65532,0,0,0,0,0,0,31,65472,0,0,0,0,0,0,31,63488,0,0,0,0,0,0,28,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	
	--944:100x9+20+20+4
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
	0,0,0,0
	);

begin
--=====================================================================================
--DHT11---------------------------
DHT11_CLK<=FD(5);	--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))操作速率
U2: DHT11_driver port Map(DHT11_CLK,DHT11_RESET,--DHT11_CLK:781250Hz(50MHz/2^6:1.28us:FD(5))操作速率,重置
						  DHT11_D_io,			--DHT11 i/o
						  DHT11_DBo,			--DHT11_driver 資料輸出
						  DHT11_RDp,			--資料讀取指標
						  DHT11_tryN,			--錯誤後嘗試幾次
						  DHT11_ok,DHT11_S,		--DHT11_driver完成作業旗標,錯誤信息						  
						  DHT11_DBoH,DHT11_DBoT,DHT11_DBoT_1,--直接輸出濕度(整數,小數固定為0值所以不輸出),溫度(整數),溫度小數1位(bit7=1為負值)
						  DHT11_DBoH1,DHT11_DBoH0,DHT11_DBoT1,DHT11_DBoT0,DHT11_DBoT_1_1,--直接輸出濕度及溫度(十位數及個位數,溫度小數1位)
						  DHT11_DBoH1_ASC,DHT11_DBoH0_ASC,DHT11_DBoT1_ASC,DHT11_DBoT0_ASC,DHT11_DBoT_1_1_ASC,--直接輸出濕度及溫度ASCII,溫度小數1位
						  H_Sound_DATA,T_Sound_DATA);--直接輸出濕度及溫度語音
--TSL2561---------------------------
--I2C2Wdriver2 介面實體
TSL2561driver:i2c2wdriver2 port map(I2CCLK=>TSL2561_CLK,			--系統時脈,系統重置
									RESET=>TSL2561_RESET,			--系統時脈,系統重置
									ID=>TSL2561_ID,					--裝置碼
									CurrentADDR=>'1',				--要求命令:(0目前位址讀取),(1指定位址讀取)
									ADDR=>TSL2561_COMMAND,			--TSL2561:COMMAND
									A2A1A0=>"001",					--ID&A2A1A0:Slave Address:0x29,0x39,0x49
									DATAin=>TSL2561_DATAin,			--資料輸入:DATA write to TSL2561
									DATAout=>TSL2561_DATAout,		--資料輸出:TSL2561 DATA read to FPGA
									RW=>TSL2561_RW,					--讀寫0:w,1:R
									RWN=>TSL2561_RWN,				--嘗試讀寫次數
									D_W_R_N=>TSL2561_D_W_R_N,		--連續讀寫次數
									D_W_R_Nok=>TSL2561_D_W_R_Nok,	--讀寫1次數旗標
									reWR=>TSL2561_reWR,				--已寫入或讀出資料
									I2Cok=>TSL2561_ok,				--TSL2561_ok 狀態
									I2CS=>TSL2561_CS,				--TSL2561_CS 狀態
									SCL=>TSL2561_SCL,				--介面IO:SCL,如有接提升電阻時可設成inout
									SDA=>TSL2561_SDA				--介面IO:SDA,有接提升電阻
									);

--SD178BMI2C---------------------------
--SD178BMI2Cdriver介面實體
SD178BMI2Cdriver1:sd178BMI2C2wdriver port map(I2CCLK=>SD178BMI2C_CLK,					--系統時脈
											  RESET=>SD178BMI2C_RESET,					--系統重置
											  ID=>SD178BMI2C_ID,						--裝置碼0100000
											  DATAin=>SD178BMI2C_DATAin,				--資料輸入
											  DATAout=>SD178BMI2C_DATAout,				--資料輸出
											  RW=>SD178BMI2C_RW,						--讀寫
											  RWN=>SD178BMI2C_RWN,						--嘗試讀寫次數
											  D_W_R_N=>SD178BMI2C_D_W_R_N,			 	--連續讀寫次數
											  D_W_R_Nok=>SD178BMI2C_D_W_R_Nok,			--讀寫1次數旗標
											  reWR=>SD178BMI2C_reWR,					--已寫入或讀出資料
											  I2Cok=>SD178BMI2C_ok,						--I2Cok
											  I2CS=>SD178BMI2C_CS,						--CS 狀態
											  SCL=>SD178BMI2C_SCL,						--介面IO:SCL,如有接提升電阻時可設成inout
											  SDA=>SD178BMI2C_SDA						--介面IO:SDA
											 );
--key board 4x4
U3: k4x4 port Map(FD(17),S_RESET,ki,ko,kn,kv,kok,koo);

--tft_lcd-------------------------------------------------------------------
st7735_spi_tft_lcd:st7735_spi_tft_lcd_4w_driver_2
			port map(st7735_CLK,st7735_RESET,	--系統時脈,系統重置
			  st7735_RES,st7735_BLS,			--介面控制:RESX,BL輸入
			  DCi,				--00:命令 01:命令參數 11:g資料
			  cmpai,			--命令_參數 輸入,水平8點image
			  cbi,				--色盤(4bit):xx01(12bit)、xx10(16bit)、xx11(18bit)
			  fcri,fcgi,fcbi,	--色系
			  bcri,bcgi,bcbi,	--色系
			  d8_1i,			--水平剩餘點數
			  --------------------------------------------------------------
			  st7735_RESX,		--介面IO:RESX輸出
			  st7735_CS,		--介面IO:CSX輸出
			  st7735_DC,		--介面IO:DCX輸出
			  st7735_SCL,		--介面IO:SCL輸出
			  st7735_SDA,		--介面IO:SDA輸出
			  st7735_BL,		--介面IO:BL輸出
			  --------------------------------------------------------------
			  st7735_reLOAD,	--載入旗標:0 可載入
			  st7735_LoadCK,	--載入時脈
			  st7735_spi_ok		--完成旗標
			);

st7735_RES<=S_RESET;

--DCmotor------------------------------------------------------------------- 
L293D: DCmotor_pwm_driver 
	port Map(FD(9),				--驅動速率
			 pwmckset,			--pwmckset:設pwm範圍0~,0:停止
			 pwmsetN,			--pwmsetN:設pwm值 ,0:停止 ,0<pwmsetN>=pwmckset:100%,1~pwmckset:pwm%
			 L293D_1A,L293D_2A,	--轉向
			 L293D_12EN			--輸出
			);

----st7735指令=========================================================================
--反相控制							--INVCTR: Display Inversion Control
st7735_IT(3)<=st7735_INVCTR;		--3 Default(03h): 0 0 0 0 0 NLA NLB NLC: 00000011
--記憶體進出入順序及顯示控制		--MADCTL (36h): Memory Data Access Control
st7735_IT(5)<=st7735_MADCTL;		--5 Default(00h): MY(0) MX(0) MV(0) ML(0) RGB(0) MH(0) - -
--色彩限定OFF(38h)／ON(39h)
st7735_IT(6)<=st7735_IDMOFF_ON;		--6 Default IDMOFF (38h)(4k,65k,262k), IDMON (39h)(only 8 color):
--不反相(20h)／反相(21h)顯示
st7735_IT(7)<=st7735_INVOFF_ON;		--7 Default INVOFF (20h): Display Inversion Off, INVON (21h): Display Inversion On
--正常(13h)／部分(12h)顯示模式
st7735_IT(8)<=st7735_NORON_PTLON;	--8 Default NORON (13h): Normal Display Mode On, PTLON (12h): Partial Display Mode On
--顯示部分範圍設定					--PTLAR
st7735_IT(11)<=CONV_STD_LOGIC_VECTOR(st7735_PSL,8);	--11 PSL7~PSL0(X"00")
st7735_IT(13)<=CONV_STD_LOGIC_VECTOR(st7735_PEL,8);	--13 PEL7~PEL0(X"A1")
--色彩深度設定 						--Interface Pixel Format:(12-bit,16-bit,18-bit)
st7735_IT(15)<=st7735_COLMOD;		--15 Default(06h):18 bit pixel format, (05h):16 bit pixel format, (03h):12 bit pixel format
----frame x範圍設定					--CASET:
st7735_IT(18)<=CONV_STD_LOGIC_VECTOR((st7735_DATA_CPOINTER_begin mod 128)+2,8);	--18 XS7~XS0(X"00")
st7735_IT(20)<=CONV_STD_LOGIC_VECTOR((st7735_DATA_CPOINTER_end mod 128)+2,8);	--20 XE7~XE0(X"83")
--frame y範圍設定					--RASET
st7735_IT(23)<=CONV_STD_LOGIC_VECTOR((st7735_DATA_RPOINTER_begin mod 160)+1,8);	--23 YS7~YS0(X"00")
st7735_IT(25)<=CONV_STD_LOGIC_VECTOR((st7735_DATA_RPOINTER_end mod 160)+1,8);	--25 YE7~YE0(X"A1")
--顯示ON/OFF設定					--27 DISPON (29h), Default DISPOFF (28h)
st7735_IT(27)<=st7735_DISPON_OFF;
--=====================================================================================
--無L293D時,運用此8pin即可(8pin排線中間線須短路，自行製作)
SD178BMI2CP_3_3V_power<=(others=>SD178BMI2CP_powerdown);

--有L293D時,如下2選1都可或接線時兩線正接或反接皆可
--SD178BMI2CP_powerdown:1:4V,0:開路
--L293D_34EN<=SD178BMI2CP_powerdown;
--L293D_3A<='1';

--SD178BMI2CP_powerdown:1:4V,0:0V
L293D_34EN<='1';
L293D_3A<=SD178BMI2CP_powerdown;--1:4V,0:0V
-----------------------------
MMx<=M710;		--M指撥開關狀態設定
-- --------------------------
E109_1_1_MainCLK<=FD(17);	--E109_1_1_Main主控器操作速率
E109_1_1_Main:process(E109_1_1_MainCLK)
variable k:integer range 0 to 31;
begin
	if S_RESET='0' then		--系統重置
		MM<=not MMx;		--虛擬指撥開關不等於實體指撥開關狀態
		D7_DB<=(0,0,0,0,0,0,0,0);	--清除顯示資料
		flash_a_g<=(others=>'0');	--off gfedcba閃爍
		flashs<=(others=>'0');		--off 小數點閃爍
		d7dot<=(others=>'0');		--off 小數點
		k:=16;						--無效鍵值
		S0on<='0';					--取消S0按鈕紀錄
		MMs<=5;						--處理結束
		Mx<=(others=>'0');			--功能執行紀錄
		SD178BMI2C_RWs<='0';		--write
		st7735_reset0<='0';			--啟動TFT_LCD首次清空
		SD178BMI2CP_reseton_delay<=0;--SD178BMI2CP_powerdown 計時歸零
	elsif rising_edge(E109_1_1_MainCLK) then

		--k4x4處理===========================
		if k/=16 then
			k:=16;
		elsif kok='1' then	--按鈕輸入
			k:=kv;
		end if;
		
		--------------------------------------------------------
		if MM/=MMx or (S0on='1' and k=0) then --實體指撥開關/=虛擬指撥開關狀態 or 測試程序停止(偵測S0on='1' and k=2)
			MM<=MMx;				--虛擬指撥開關等於實體指撥開關狀態
			S0on<='0';				--取消按鈕紀錄
			-------------------------------------------
			DHT11_RESET<='0';		--DHT11_driver控制旗標
			-------------------------------------------
			TSL2561P_reset<='0';	--TSL2561_P控制旗標 TSL2561_P off
			-------------------------------------------
			SD178BMI2CP_reset<='0'; --SD178BMI2CP off
			SD178BMI2CP_reseton<='0';--執行"硬體reset"
			SD178BMI2CP_powerdown<='1';--電源重啟:off
			SD178BMI2C_sound(0 to 1)<=(X"01",X"80");--V2版(X"01",X"80"):會當機(死當)
			--(X"00",X"00")硬體reset or (X"00",X"01")nop or 任一立即執行命令:如(X"01",X"80")都ok;但V2版只有(X"01",X"80":會當機)已轉成"硬體reset"操作(防當機)
			SD178BMI2C_P_end_t_onoff<='0';	--off 是否啟動終止延遲計時
			SD178BMI2C_P_end_t_set<=0;		--0,終止延遲計時次數(1:約1.004ms)
			-------------------------------------------
			st7735_P_RESET<='0';			--st7735_P off
			st7735_BLS<='1';				--背光on
			st7735_DATA_C_INC<=16;			--1~16
			st7735_COLMOD<=X"05";			--15 Default(06h)(18-bit/pixel)=R(6bit)G(6bit)B(6bit):(X"06"18-bit)(X"05"16-bit)(X"03"12-bit);
			st7735_INVCTR<=X"03";			--3 Default(03h): 0 0 0 0 0 NLA NLB NLC: 00000011
			st7735_MADCTL<=X"C0";			--4 Default(00h):MY(0) MX(0) MV(0) ML(0) RGB(0) MH(0) - -
			st7735_IDMOFF_ON<=X"38";		--6 Default IDMOFF (38h)(4k,65k,262k), IDMON (39h)(only 8 color)
			st7735_INVOFF_ON<=X"20";		--7 Default INVOFF (20h): Display Inversion Off, INVON (21h): Display Inversion On
			st7735_NORON_PTLON<=X"13";		--8 Default NORON (13h): Normal Display Mode On, PTLON (12h): Partial Display Mode On
			st7735_DISPON_OFF<=X"29";		--27 DISPON (29h), Default DISPOFF (28h)
			st7735_PSL<=0;					--列起點
			st7735_PEL<=161;				--列終點
			st7735_DATA_CPOINTER_begin<=0;	--行起點
			st7735_DATA_RPOINTER_begin<=0;	--列起點
			st7735_DATA_CPOINTER_end<=127;	--行終點 128:0~127
			st7735_DATA_RPOINTER_end<=159;	--列終點 160:0~159
			if st7735_reset0='0' then
				st7735_COM_POINTERs<=0;		--tft lcd命令指標
				SD178BMI2CP_powerdown<='0';--電源重啟:on
			else
				st7735_COM_POINTERs<=16;	--tft lcd命令指標
			end if;
			st7735_time_Dn<=0;				--完成後延遲時間設定
			B1_COLORi<=0;					--1選色 黑
			B0_COLORi<=7;					--0選色 白
			monoC<=0;						--單色操作
			isword<=false;					--圖形或字型:圖形
			remove_leading_0<='0';			--去前導零off
			word_w<=20;						--字寬
			gdata0<=(others=>'0');			--單色圖樣	
			cbis<="0010";					--色盤:單色16bit
			st7735_ch<="0000";				--ch="0000"
		elsif SD178BMI2CP_powerdown='0' or SD178BMI2CP_reseton_delay/=0 then
			SD178BMI2CP_reseton_delay<=SD178BMI2CP_reseton_delay-1;
			SD178BMI2CP_reset<='0'; --SD178BMI2CP off
			if SD178BMI2CP_reseton_delay=0 then
				SD178BMI2CP_reseton<='0';--SD178BMI2C 硬體reset
				SD178BMI2CP_reseton_delay<=80;
			end if;
			if SD178BMI2CP_reseton_delay=70 then
				SD178BMI2CP_powerdown<='1';
			end if;
			if SD178BMI2CP_reseton_delay=45 then
				SD178BMI2CP_reseton<='1';
			end if;
			
		elsif SD178BMI2CP_reseton='0' then	--未啟動SD178BMI2CP執行硬體reset
			SD178BMI2CP_reseton_delay<=60;

		elsif st7735_reset0='0' then	--TFT_LCD首次清空
			if st7735_P_ok='1' then
				st7735_reset0<='1';
				st7735_P_RESET<='0';
			else
				gdata0<=(others=>'0');	--單色圖樣(全白)
				st7735_P_RESET<='1';
			end if;
 		else
			--s2(停止鍵)再按下之後,按S1(重置鍵)回到該功能初始設定狀態之處理
			if (Mx(conv_integer(MMx))='1' and k=1 and S0on='0') or MMs=6 then
				if MMs=5 then
					st7735_COM_POINTERs<=16;		--tft lcd命令指標:16 CASET(2Ah): Column Address Set
					st7735_P_RESET<='1';
					D7_DB<=(others=>0);		--顯示預設值00000000
					flash_a_g<=(others=>'0');--off gfedcba閃爍
					flashs<=(others=>'0');	--off--小數點無閃爍
					d7dot<=(others=>'0');	--off--小數點
					case MMx is
						when "00"=>
							Mx(0)<='0';
						when "01"=>
--							D7_DB<=(others=>0);		--顯示預設值00000000
--							flash_a_g<=(others=>'0');--off gfedcba閃爍
--							flashs<=(others=>'0');	--off--小數點無閃爍
--							d7dot<=(others=>'0');	--off--小數點
							Mx(1)<='0';
						when "10"=>
							Mx(2)<='0';
						when others=>
							gdata0<=(others=>'1');	--單色圖樣(全黑)
							Mx(3)<='0';
					end case;
					MMs<=6;					--繼續下一步
				elsif st7735_P_ok='1' then
					MMs<=5;					--處理結束
					st7735_P_RESET<='0';
				end if;
			else
				---------------------------------------------------------------------------------------
				--00 or 11 LCD秀
				if (MMx=0 or MMx=3)and S0on='1' and times1<18 then
					if st7735_P_ok='1' then
						st7735_COM_POINTERs<=21;		--tft lcd命令指標:21 RASET(2Bh): Row Address Set
						times1<=times1-1;	--下一步
						if times1=1 then
							times1<=17;		--顯示重來
						end if;
						if times1>9 then--17..10白<->黑 17 16 15 14 13 12 11 10
							st7735_ch<="0000";					--ch0
							if times1 mod 2=1 then --17 15 13 11
								st7735_DATA_RPOINTER_begin<=0;	--列起點
								st7735_DATA_RPOINTER_end<=79;	--列終點
								st7735_time_Dn<=0;				--完成後延遲時間設定0s
							else --16 14 12 10
								st7735_DATA_RPOINTER_begin<=80;	--列起點
								st7735_DATA_RPOINTER_end<=159;	--列終點
								st7735_time_Dn<=50000000;		--完成後延遲時間設定0.5s
								B0_COLORi<=7-B0_COLORi;			--0選色:白7/黑0(白<->黑)
							end if;
							if times1=17 then	--顏色初值預設
								B0_COLORi<=7;	--0選色:白7
								B1_COLORi<=0;	--0選色:黑0
							end if;
						elsif times1 <= 3 then -- 9..1
							st7735_ch<="0001";				--ch1
							st7735_time_Dn<=50000000;		--完成後延遲時間設定1s
							st7735_DATA_RPOINTER_begin<=0;	--列起點
							st7735_DATA_RPOINTER_end<=159;	--列終點
							B0_COLORi<=7;					--0選色:白7
							if times1<4 then
								B1_COLORi<= 4 - times1;			--1選色:B3,G2,R1
							end if;
							beFriendC_P<=1280* (4 - times1) +80;	--大字:123456789
						end if;
						st7735_P_RESET<='0';	--off
					else
						st7735_P_RESET<='1';	--on
					end if;
				end if;
			---------------------------------------------------------------------------------------
	
				case MMx is
					--00--TFT_LCD test---------------------------------
					when "00" =>	--由按s0起動 TFT_LCD test
						if S0on='0' then
							st7735_COM_POINTERs<=16;	--tft lcd命令指標:16 CASET(2Ah): Column Address Set
							if k=0 then	--偵測k=0 start
								S0on<='1';	--紀錄S0on
								Mx(0)<='1';	--功能執行紀錄:恢復旗標
								D7_DB<=(others=>0);		--顯示預設值00000000
								d7dot<=(others=>'0');	--off--小數點
								times1<=18;				--顯示步驟預設
							end if;
						elsif k=1 then	--偵測k=1重置
							st7735_COM_POINTERs<=16;		--tft lcd命令指標:16 CASET(2Ah): Column Address Set
							st7735_DATA_CPOINTER_begin<=0;	--行起點
							st7735_DATA_CPOINTER_end<=127;	--行終點 128:0~127
							st7735_DATA_RPOINTER_begin<=0;	--列起點
							st7735_DATA_RPOINTER_end<=159;	--列終點 160:0~159
							times1<=18;						--顯示重來
							st7735_ch<="0000";				--ch0
							st7735_time_Dn<=0;				--完成後延遲時間設定0s
							st7735_P_RESET<='0';			--off
--						elsif st7735_P_ok='1' then
--							st7735_COM_POINTERs<=21;		--tft lcd命令指標:21 RASET(2Bh): Row Address Set
--							times1<=times1-1;	--下一步
--							if times1=1 then
--								times1<=17;		--顯示重來
--							end if;
--							if times1>9 then--17..10白<->黑
--								st7735_ch<="0000";					--ch0
--								if times1 mod 2=1 then
--									st7735_DATA_RPOINTER_begin<=0;	--列起點
--									st7735_DATA_RPOINTER_end<=79;	--列終點
--									st7735_time_Dn<=0;				--完成後延遲時間設定0s
--								else
--									st7735_DATA_RPOINTER_begin<=80;	--列起點
--									st7735_DATA_RPOINTER_end<=159;	--列終點
--									st7735_time_Dn<=50000000;		--完成後延遲時間設定0.5s
--									B0_COLORi<=7-B0_COLORi;			--0選色:白7/黑0(白<->黑)
--								end if;
--								if times1=17 then	--顏色初值預設
--									B0_COLORi<=7;	--0選色:白7
--									B1_COLORi<=0;	--0選色:黑0
--								end if;
--							else	--9..1
--								st7735_ch<="0001";				--ch1
--								st7735_time_Dn<=50000000;		--完成後延遲時間設定1s
--								st7735_DATA_RPOINTER_begin<=0;	--列起點
--								st7735_DATA_RPOINTER_end<=159;	--列終點
--								B0_COLORi<=7;					--0選色:白7
--								if times1<4 then
--									B1_COLORi<=times1;			--1選色:B3,G2,R1
--								end if;
--								beFriendC_P<=1280*times1+80;		--大字:123456789
--							end if;
--							st7735_P_RESET<='0';	--off
--						else
--							st7735_P_RESET<='1';	--on
						elsif times1=18 then
							st7735_P_RESET<='1';	--清空LCD
							times1<=17;
						end if;

					--01--SD178BMI2C 音量、聲道測試---------------------------------
					when "01" =>	--由按S0起動
						if S0on='0' then
							st7735_COM_POINTERs<=16;	--tft lcd命令指標:16 CASET(2Ah): Column Address Set
							if k=0 then	--偵測k=0 start
								S0on<='1';	--紀錄S0on
								Mx(1)<='1';	--功能執行紀錄:恢復旗標
								F12<=0;		--預設音量功能
								F1<=3;		--預設音量
								F2<=1;		--預設聲道
													 --0  1  2  3  4  5  6  7  8  9
								Sound86<=3;	--預設音量 00 87 96 A5 B4 C3 D2 E1 F0 FF 每階15
								Sound8B<=1;	--預設聲道
							end if;
						elsif k=1 then	--偵測k=1重置
							F12<=0;		--預設音量功能
							F1<=3;		--預設音量
							F2<=1;		--預設聲道
												 --0  1  2  3  4  5  6  7  8  9
							Sound86<=3;	--預設音量 00 87 96 A5 B4 C3 D2 E1 F0 FF 每階15
							Sound8B<=1;	--預設聲道
							SD178BMI2CP_powerdown<='0';	--電源重啟:on(語音模組重啟防當機)
							st7735_P_RESET<='0';		--off
						else
							st7735_P_RESET<='1';
							if SD178BMI2CP_ok='1' then
								if F12=0 then
									D7_DB<=(F1,0,13,0,15,16,1,11);	--顯示預設值F1.VOL03
									d7dot<="11111011";				--off--小數點
									if k=4 then		--up不可循環設計
										if F1/=9 then
											F1<=F1+1;
										end if;
									elsif k=5 then	--down不可循環設計
										if F1/=0 then
											F1<=F1-1;
										end if;
									end if;
								else
									if F2=1 then
										D7_DB<=(7,12,6,1,14,16,2,11);	--顯示預設值F2.RIGH(T.)
										d7dot<="01111011";				--off--小數點
									elsif F2=2 then
										D7_DB<=(16,7,11,10,13,16,2,11);	--顯示預設值F2.LEF(T.).
										d7dot<="00111011";				--off--小數點
									else
										D7_DB<=(16,12,7,0,8,16,2,11);	--顯示預設值(F.)2.BOTH.
										d7dot<="01111010";				--off--小數點
									end if;
									if k=4 then		--up可循環設計
										if F2=1 then
											F2<=3;
										else
											F2<=F2-1;
										end if;
									elsif k=5 then	--down可循環設計
										if F2=3 then
											F2<=1;
										else
											F2<=F2+1;
										end if;
									end if;
								end if;
								if k=2 then		--切換功能
									F12<=1-F12;	--0/1
								elsif k=6 then	--設定功能
									if F12=0 then
										Sound86<=F1;
									else
										-- {{ by myself start }}
										if F2=1 then
											Sound8B<=2;
										elsif F2=2 then
											Sound8B<=1;
										else
											Sound8B<=3;
										end if;
										-- {{ by myself end }}
										-- Sound8B<=F2;
									end if;
									SD178BMI2CP_reset<='0';	--on
								end if;								
							else
								SD178BMI2CP_reset<='1';	--on
								SD178BMI2C_sound(0 to 11)<=(X"0B",X"8F",X"02",--Skip 提前結束正執行的87H或88H指令，跳至下一指令
															X"86",Sound86_VOL(Sound86),X"8B",Sound8B_R_L(Sound8B),--86:音量 5->D7 8B:RL聲道設定
															X"88",X"23",X"38",X"00",X"00");--選曲0~9:9008~9017(X"2330"~X"2339")無限次
							end if;
						end if;

					--10--TSL2561 & DHT11 test---------------------------------
					when "10" =>	--由按0起動
						if S0on='0' then
							st7735_COM_POINTERs<=16;	--tft lcd命令指標:16 CASET(2Ah): Column Address Set
							if k=0 then	--偵測k=0 start
								S0on<='1';	--紀錄S0on
								Mx(2)<='1';	--功能執行紀錄:恢復旗標
								D7_DB<=(others=>0);		--顯示預設值00000000
								d7dot<=(others=>'0');	--off--小數點
								remove_leading_0<='1';	--去前導零on
							end if;
							times<=100;
						elsif k=1 then	--偵測k=1重置
							st7735_COM_POINTERs<=16;		--tft lcd命令指標:16 CASET(2Ah): Column Address Set
							st7735_DATA_CPOINTER_begin<=0;	--行起點
							st7735_DATA_CPOINTER_end<=127;	--行終點 128:0~127
							st7735_DATA_RPOINTER_begin<=0;	--列起點
							st7735_DATA_RPOINTER_end<=159;	--列終點 160:0~159
							gdata0<=(others=>'0');			--單色圖樣(全白)
							st7735_ch<="0000";				--ch="0000"
							isword<=false;					--圖形或字型:字型
							st7735_P_RESET<='0';
							DHT11_RESET<='0';		--off
							TSL2561P_reset<='0';	--off
							times<=100;
						elsif st7735_P_ok='1' then
							if TSL2561P_reset='0' or DHT11_RESET='0' then	--尚未啟動讀取感測器數據
								TSL2561P_reset<='1';	--起動 TSL2561_P
								DHT11_RESET<='1';		--起動 DHT11_driver
							elsif TSL2561P_ok='1' and DHT11_ok='1' then		--已完成讀取感測器數據
								times<=times-1;	--計時
								if times=0 then
									DHT11_RESET<='0';		--off
									TSL2561P_reset<='0';	--off
									times<=100;
--								elsif DHT11_S='1' then	--資料讀取失敗
--									null;				
								else
									st7735_ch<="0010";		--ch="0010"
									B1_COLORi<=0;			--1選色(黑)
									isword<=true;			--圖形或字型:字型
									word_w<=20;				--字寬
									beFriendC_P<=0;
									if times=100 then--亮度
										st7735_DATA_CPOINTER_begin<=0;	--行起點
										st7735_DATA_CPOINTER_end<=99;	--行終點
										st7735_DATA_RPOINTER_begin<=0;	--列起點
										st7735_DATA_RPOINTER_end<=39;	--列終點
										st7735_P_RESET<='0';
										if M70s(4)(2)='1' then
											st7735_DATA<=(LUX(3),LUX(2),LUX(1),10,LUX(0));
										else
											st7735_DATA<=(2,3,3,1,0);
											st7735_DATA_CPOINTER_end<=127;	--行終點
											word_w<=32;			--字寬
											B1_COLORi<=1;		--1選色(紅)
											beFriendC_P<=800;
										end if;
										
									elsif times=99 then--溫度
										st7735_DATA<=(0,DHT11_DBoT1,DHT11_DBoT0,10,DHT11_DBoT_1_1);
										st7735_DATA_CPOINTER_begin<=0;	--行起點
										st7735_DATA_CPOINTER_end<=99;	--行終點
										st7735_DATA_RPOINTER_begin<=60;	--列起點
										st7735_DATA_RPOINTER_end<=99;	--列終點
										st7735_P_RESET<='0';
										if M70s(3)(2)='1' then
											st7735_DATA<=(0,DHT11_DBoT1,DHT11_DBoT0,10,DHT11_DBoT_1_1);
										else
											st7735_DATA<=(2,3,3,1,0);
											st7735_DATA_CPOINTER_end<=127;	--行終點
											word_w<=32;			--字寬
											B1_COLORi<=2;		--1選色(綠)
											beFriendC_P<=800;
										end if;

									elsif times=98 then--濕度
										st7735_DATA<=(0,DHT11_DBoH1,DHT11_DBoH0,10,0);
										st7735_DATA_CPOINTER_begin<=0;	--行起點
										st7735_DATA_CPOINTER_end<=99;	--行終點
										st7735_DATA_RPOINTER_begin<=120;--列起點
										st7735_DATA_RPOINTER_end<=159;	--列終點
										st7735_P_RESET<='0';
										if M70s(2)(2)='1' then
											st7735_DATA<=(0,DHT11_DBoH1,DHT11_DBoH0,10,0);
										else
											st7735_DATA<=(2,3,3,1,0);
											st7735_DATA_CPOINTER_end<=127;	--行終點
											word_w<=32;			--字寬
											B1_COLORi<=3;		--1選色(藍)
											beFriendC_P<=800;
										end if;

									elsif times=97 then--亮度Lux.1120
										st7735_DATA_CPOINTER_begin<=100;--行起點
										st7735_DATA_CPOINTER_end<=127;	--行終點
										if M70s(4)(2)='1' then
											beFriendC_P<=1120;
											st7735_DATA_RPOINTER_begin<=0;	--列起點
											st7735_DATA_RPOINTER_end<=39;	--列終點
											st7735_ch<="0001";	--ch="0001"
											B1_COLORi<=1;		--1選色(紅)
											isword<=false;			--圖形或字型:圖形
											st7735_P_RESET<='0';
										end if;

									elsif times=96 then--溫度℃1200
										if M70s(3)(2)='1' then
											beFriendC_P<=1200;
											st7735_DATA_RPOINTER_begin<=60;	--列起點
											st7735_DATA_RPOINTER_end<=99;	--列終點
											st7735_ch<="0001";	--ch="0001"
											B1_COLORi<=2;		--1選色(綠)
											isword<=false;			--圖形或字型:圖形
											st7735_P_RESET<='0';
										end if;

									elsif times=95 then--濕度%1280
										if M70s(2)(2)='1' then
											beFriendC_P<=1280;
											st7735_DATA_RPOINTER_begin<=120;	--列起點
											st7735_DATA_RPOINTER_end<=159;	--列終點
											st7735_ch<="0001";	--ch="0001"
											B1_COLORi<=3;		--1選色(藍)
											isword<=false;			--圖形或字型:圖形
											st7735_P_RESET<='0';
										end if;
									
									end if;
								end if;
							end if;
						else
							st7735_P_RESET<='1';
						end if;

					--11--SD178BMI2C 語音播放 test---------------------------------
					when "11" =>
						if S0on='0' then
							st7735_COM_POINTERs<=16;	--tft lcd命令指標:16 CASET(2Ah): Column Address Set
							if k=0 then	--偵測k=0 start
								S0on<='1';	--紀錄S0on
								Mx(3)<='1';	--功能執行紀錄:恢復旗標
								soundn<=0;
								D7_DB<=(others=>0);		--顯示預設值00000000
								d7dot<=(others=>'0');	--off--小數點
								times1<=18;				--LCD顯示重來
							end if;
						elsif k=1 then	--偵測k=1重置
							soundn<=0;
							SD178BMI2C_sound(0 to 1)<=(X"00",X"00");--(X"00",X"00")硬體reset
							SD178BMI2CP_reset<='0';							
							SD178BMI2C_P_end_t_set<=0;	--0,終止延遲計時次數(1:約1.004ms)
							st7735_ch<="0000";			--ch0
							times1<=18;					--LCD顯示重來
							st7735_P_RESET<='0';		--off
						else
							if times1=18 then
								st7735_P_RESET<='1';	--清空LCD
								times1<=17;
							end if;
							if SD178BMI2CP_ok='1' then
								SD178BMI2CP_reset<='0';	--off
								SD178BMI2C_P_end_t_onoff<='1';	--off 是否啟動終止延遲計時
								SD178BMI2C_P_end_t_set<=1000;	--0,終止延遲計時次數(1:約1.004ms)
								soundn<=soundn+1;
								case soundn is
									when 0=>
									--撥放”系統開機”
									SD178BMI2C_sound(0 to 21)<=(X"19",X"86",X"D7",X"8B",X"07",--86:音量 5->D7 8B:RL聲道設定 
																-- X"BC",X"BD",X"A9",X"F1",--播放
																X"87",X"00",X"00",X"03",X"E8",--delay 1s
																X"A8",X"74",X"B2",X"CE",X"B6",X"7D",X"BE",X"F7",--系統開機
																X"8A",X"06",X"8A",X"07");--等待撥音結束

									when 1=>
									--播放”撥放右左或雙聲道”
									SD178BMI2C_sound(0 to 24)<=(X"20",X"86",X"D7",X"8B",X"07",--86:音量 5->D7 8B:RL聲道設定 
																-- X"BC",X"BD",X"A9",X"F1",--播放
																X"87",X"00",X"00",X"03",X"E8",--delay 1s
																-- X"A5",X"6B",--右
																X"BC", X"C6", X"A6", X"72", X"B4", X"FA", X"B8", X"D5", -- 系統測試
																X"87",X"00",X"00",X"01",X"f4",--delay 0.5s
																-- X"A5",X"AA",X"A9",X"CE",X"C2",X"F9",X"C1",X"6E",X"B9",X"44",--左或雙聲道
																X"8A",X"06");--等待撥音結束
									when 2=>
									--播放”感測器的數值與設定”
									SD178BMI2C_sound(0 to 35)<=(X"23",X"86",X"D7",X"8B",X"07",--86:音量 5->D7 8B:RL聲道設定 
																X"BC",X"BD",X"A9",X"F1",--播放
																X"87",X"00",X"00",X"03",X"E8",--delay 1s
																X"B7",X"50",X"B4",X"FA",X"BE",X"B9",X"AA",X"BA",X"BC",X"C6",X"AD",X"C8",X"BB",X"50",X"B3",X"5D",X"A9",X"77",--感測器的數值與設定
																X"8A",X"06",X"8A",X"07");--等待撥音結束
									when others=>
									--播放”再測試一次”
									SD178BMI2C_sound(0 to 27)<=(X"1B",X"86",X"D7",X"8B",X"07",--86:音量 5->D7 8B:RL聲道設定 
																X"BC",X"BD",X"A9",X"F1",--播放
																X"87",X"00",X"00",X"03",X"E8",--delay 1s																
																X"A6",X"41",X"B4",X"FA",X"B8",X"D5",X"A4",X"40",X"A6",X"B8",--再測試一次
																X"8A",X"06",X"8A",X"07");--等待撥音結束
									soundn<=0;
								end case;
							else
								SD178BMI2CP_reset<='1';	--on
							end if;
						end if;

------------------------------------------------------------------------------------------------------------------------
					when others =>	
						null;
				end case;
			end if;
		end if;
	end if;
end process E109_1_1_Main;

--=====================================================================================
--七段顯示器---------------------------------------------------
--8位數掃瞄器
scan_P:process(FD(14),S_RESET)
begin
	if S_RESET='0' then
		scanP<=0;		--位數取值指標
		SCANo<="00000000";	--掃瞄信號
	elsif rising_edge(FD(14)) then
		scanP<=scanP+1;
		SCANo<=SCANo(6 downto 0)&SCANo(7);
		if scanP=7 then
			scanP<=0;
			SCANo<="11111110";--掃瞄信號
		end if;
	end if;
end process scan_P;

--BCD碼解共陽極七段顯示碼pgfedcba:d7dot(scanP)=1有小數點 ,flashs(scanP)=1小數點閃爍
flash_a_gs<="1111111" when (flash_a_g(scanP) and FD(23))='1' else "0000000";--gfedcba閃爍
D7LED<=(not d7dot(scanP)or(d7dot(scanP)and flashs(scanP)and FD(23)))
	 & (Disp7(D7_DB(scanP))or flash_a_gs);
D7LED2<=(not d7dot(scanP)or(d7dot(scanP)and flashs(scanP)and FD(23)))
	 & (Disp7(D7_DB(scanP))or flash_a_gs);
--=====================================================================================
--tft lcd顯示器
--頁顯示資料解碼
--去前導零xxx.x
st7735_x0<=0 when st7735_DATA(0)>0  or remove_leading_0='0' else
		   1 when st7735_DATA(1)>0 else
		   2;

--查字:isword=true
gdata2<=CONV_STD_LOGIC_VECTOR(beFriend(beFriendC_P
									   +st7735_DATA(st7735_x/W_w_b)*W_w_b*(st7735_DATA_RPOINTER_end-st7735_DATA_RPOINTER_begin+1)
									   +(st7735_x mod W_w_b)
									   +st7735_y*W_w_b)
							  ,16)  
		when st7735_x/W_w_b>=st7735_x0 else (others=>'0');

--查圖:isword=false
gdata1<=CONV_STD_LOGIC_VECTOR(beFriend(beFriendC_P+st7735_xinc1),16);
--tft lcd顯示器================
--單色圖
with st7735_ch select
gdata<=gdata0	 when "0000",
	   gdata1 	 when "0001",
	   gdata2 	 when "0010",
	   gdata3 	 when "0011",
	   gdata4 	 when "0100",
	   gdata5 	 when "0101",
	   gdata6 	 when "0110",
	   gdata7 	 when "0111",
	   "1111111111111111"when "1000",
	   gdata9 	 when "1001",
	   gdata10 	 when others;

--色盤-------------------------
cbi<=cbis;

--單色圖1配色 或 彩色圖色------
fcri<=st7735_8baseCOLOR(B1_COLORi)(0) when monoC=0 else fc2(0);
fcgi<=st7735_8baseCOLOR(B1_COLORi)(1) when monoC=0 else fc2(1);
fcbi<=st7735_8baseCOLOR(B1_COLORi)(2) when monoC=0 else fc2(2);
--單色圖0配色---------------
bcri<=st7735_8baseCOLOR(B0_COLORi)(0) when monoC=0 else bc2(0);
bcgi<=st7735_8baseCOLOR(B0_COLORi)(1) when monoC=0 else bc2(0);
bcbi<=st7735_8baseCOLOR(B0_COLORi)(2) when monoC=0 else bc2(0);

--==========================
--單色圖水平剩餘點數解碼:st7735_DATA_C_INC:1~16
d8_1i<=(word_w mod 16)		when isword and (word_w mod 16)/=0 and (st7735_x mod W_w_b)=W_w_b-1 else
		st7735_DATA_C_INC	when st7735_DATA_CPOINTER+st7735_DATA_C_INC-1<=st7735_DATA_CPOINTER_end
							else st7735_DATA_CPOINTER_end-st7735_DATA_CPOINTER+1;
--字型word							
W_w_b<=word_w/16 when (word_w mod 16)=0 else (word_w/16)+1;

-------命令-----------------------------------------------單色圖
cmpai<="00000000"&st7735_IT(st7735_COM_POINTER) when DCi(1)='0' else gdata;

-------命令參數解碼---------------------------------------------------
with st7735_IT(st7735_COM_POINTER) select	--only write command
st7735_COM_PN0<=1	when X"26", --GAMSET
				4	when X"2A", --CASET
				4	when X"2B", --RASET
				31	when X"2C", --SW:=false;--RAMWR 準備傳送顯示資料
				4	when X"30", --PTLAR
				1	when X"36", --MADCTL
				1	when X"3A", --COLMOD
				3	when X"B1", --FRMCTR1
				3	when X"B2", --FRMCTR2
				6	when X"B3", --FRMCTR3
				1	when X"B4", --INVCTR
				2	when X"B6", --DISSET5
				2	when X"C0", --PWCTR1
				1	when X"C1", --PWCTR2
				4	when X"C2", --PWCTR3
				4	when X"C3", --PWCTR4
				2	when X"C4", --PWCTR5
				2	when X"C5", --VMCTR1
				1	when X"C7", --VMOFCTR
				16	when X"E0", --GAMCTRP1
				16	when X"E1", --GAMCTRN1
				2	when X"FC", --PWCTR6
				3	when X"FF", --VCOM4L
				0	when others;--others command

--------------------------------------------------------------
st7735_CLK<=SCLK;			--st7735操作速率
st7735_P_CLK<=SCLK;			--st7735_P操作速率
st7735_P:process(st7735_P_CLK,st7735_P_RESET)
	variable SW:Boolean;	--狀態控制旗標
	variable SWok:std_logic;--完成控制旗標
	variable td:integer range 0 to 100000000;
begin
	if st7735_P_RESET='0' then
		st7735_RESET<='0';		--st7735_spi_tft_lcd_4w_driver重置
		st7735_COM_POINTER<=st7735_COM_POINTERs;--命令起點
		st7735_LoadCK<='0';		--Load CK
		st7735_COM_PN<=st7735_COM_PN0;
		SW:=true;				--載入狀態旗標
		if st7735_COM_PN0=31 then
			SW:=false;			--載入狀態旗標
		end if;
		st7735_x<=0;			--行x POINTER
		st7735_y<=0;			--列y POINTER
		st7735_xincN<=0;		--行x incN POINTER
		st7735_xinc1<=0;		--列x inc 1... POINTER
		st7735_P_ok<='0';		--st7735_P 完成指標
		SWok:='0';
		DCi<="00";				--DC--命令參數解碼
		td:=st7735_time_Dn;		--完成後延遲時間<=2S
	elsif rising_edge(st7735_P_CLK) then
		st7735_LoadCK<='0';
		if SWok='1' then
			if td=0 then
				st7735_P_ok<='1';	--結束
			else
				td:=td-1;
			end if;
		elsif st7735_RESET='0' then
			st7735_RESET<='1';		--啟動 st7735_spi_tft_lcd_4w_driver
			st7735_DATA_CPOINTER<=st7735_DATA_CPOINTER_begin;--行起點
			st7735_DATA_RPOINTER<=st7735_DATA_RPOINTER_begin;--列起點
		elsif st7735_COM_POINTER<st7735_IT'length and st7735_COM_PN/=31 then	--傳送命令
			if st7735_COM_PN=0 then
				DCi<="00";	--DC--命令參數解碼
			else
				DCi<="01";	--DC--命令參數解碼
			end if;
			if SW=true then
				st7735_COM_POINTER<=st7735_COM_POINTER+1;
				SW:=false;
			elsif st7735_reLOAD='0' then--載入
				st7735_LoadCK<='1';
				SW:=true;
				if st7735_COM_PN/=0 then
					st7735_COM_PN<=st7735_COM_PN-1;
				else	--命令參數解碼
					st7735_COM_PN<=st7735_COM_PN0;
					if st7735_COM_PN0=31 then	--RAMWR 準備傳送顯示資料
						SW:=false;				--載入狀態旗標
					end if;
				end if;
			end if;
		elsif st7735_COM_PN/=31 then	--只下指令
			SWok:=st7735_spi_ok;	--等待結束
		elsif st7735_DATA_RPOINTER<=st7735_DATA_RPOINTER_end then	--傳送顯示資料(畫面更新)
			DCi<="11";	--DC--命令參數解碼 顯示資料
			if SW then
				if isword and (word_w mod 16)/=0 and (st7735_x mod W_w_b)=W_w_b-1 then
					st7735_DATA_CPOINTER<=st7735_DATA_CPOINTER+(word_w mod 16);			--下一行或段
					st7735_xincN<=st7735_xincN+(word_w mod 16);
				else					
					st7735_DATA_CPOINTER<=st7735_DATA_CPOINTER+st7735_DATA_C_INC;			--下一行或段
					st7735_xincN<=st7735_xincN+st7735_DATA_C_INC;
				end if;
				st7735_x<=st7735_x+1;
				st7735_xinc1<=st7735_xinc1+1;
				if st7735_DATA_CPOINTER+st7735_DATA_C_INC>st7735_DATA_CPOINTER_end then	--資料換頁
					st7735_DATA_CPOINTER<=st7735_DATA_CPOINTER_begin;
					st7735_xincN<=0;
					st7735_x<=0;
					st7735_DATA_RPOINTER<=st7735_DATA_RPOINTER+1;--資料換頁 下一ROW
					st7735_y<=st7735_y+1;
				end if;
				SW:=false;				--載入狀態旗標
			elsif st7735_reLOAD='0' and DCi="11" then
				st7735_LoadCK<='1';
				SW:=true;				--載入狀態旗標
			end if;
		else
			SWok:=st7735_spi_ok;	--等待結束
		end if;
	end if;
end process st7735_P;

--=====================================================================================
--TSL2561--------------------------------------
TSL2561_CLK<=FD(8);	--I2C時脈
TSL2561_P:process(FD(9))
variable TSL2561P_case:integer range 0 to 7;
variable LST_time:integer range 0 to 63;
begin
	if  TSL2561P_reset='0' then
		TSL2561P_case:=0;
		TSL2561P_ok<='0';		--TSL2561_P 完成指標
		TSL2561_RESET<='0';		--i2c2wdriver2重置
		TSL2561_reWR<='0';		--繼續
		TSL2561_COMMAND<="11000000";	--clear
		TSL2561_DATAin<=(others=>'0');	--power down
		TSL2561_RW<='0';		--write
		TSL2561_D_W_R_N<=1;		--單獨操作1筆
		LST_time:=31;			--delay
		TSL2561_DP<=0;
	elsif rising_edge(FD(9)) then
		if TSL2561P_ok='0' then
			if TSL2561_reWR='1' then
				TSL2561_reWR<='0';		--page作業:繼續
			elsif TSL2561_RESET='0' then
				TSL2561_RESET<='1';		--啟動i2c2wdriver2
			elsif TSL2561_ok='1' then	--完成
				case TSL2561P_case is
					when 0=>	--clera INT and power off -> clera INT and power up
						LST_time:=LST_time-1;
						if LST_time=0 then
							TSL2561_DATAin<=X"03";	--power on
							TSL2561_RESET<='0';		--i2c2wdriver2重置
							TSL2561P_case:=1;		--next step
						end if;

					when 1=>	--set INT:clera INT and level interrupt enable
							TSL2561_COMMAND<="11000110";	--clear and 06
							TSL2561_DATAin<=X"10";			--level interrupt enable
							TSL2561_RESET<='0';				--i2c2wdriver2重置
							TSL2561P_case:=2;				--next step

					when 2=>	--read DATA0LOW,DATA0HIGH,DATA1LOW,DATA1HIGH
						if TSL2561_INT='0' then
							TSL2561_COMMAND<="10001100";	--DATA0LOW:C
							TSL2561_RW<='1';				--read
							TSL2561_D_W_R_N<=4;				--操作4筆
							TSL2561_RESET<='0';				--i2c2wdriver2重置
							TSL2561P_case:=3;				--next step
						end if;

					when 3=>	--clera INT and power off
						TSL2561_DATA01(TSL2561_DP)<=TSL2561_DATAout;--輸出資料
						TSL2561_COMMAND<="11000000";	--clear INT
						TSL2561_DATAin<=(others=>'0');	--power down
						TSL2561_RW<='0';				--write
						TSL2561_D_W_R_N<=1;				--操作1筆
						TSL2561_RESET<='0';				--i2c2wdriver2重置
						TSL2561P_case:=4;				--next step

					when others=>	--TSL2561_P 完成
						TSL2561P_ok<='1';		--TSL2561_P 完成指標
						TSL2561_RESET<='0';		--i2c2wdriver2重置

				end case;
			elsif TSL2561_D_W_R_Nok='1' then		--page作業通知
				TSL2561_DATA01(TSL2561_DP)<=TSL2561_DATAout;--輸出資料
				TSL2561_DP<=TSL2561_DP+1;			--下一筆
				TSL2561_reWR<='1';					--回收到
			end if;
		end if;
	end if;
end process TSL2561_P;

---------------------------------------------------------------------------------------------------
--計算TSL2561照度值
--iGain 0:=1X 1:16X ,Tint 0:=13.7ms, 1:101ms, 2:402ms ,iType 0:T,FN,CL 1:CS
--default
--iGain:0			,Tint:2							  ,iType:0
CH0<=conv_integer(TSL2561_DATA01(1)&TSL2561_DATA01(0));	--16bit
CH1<=conv_integer(TSL2561_DATA01(3)&TSL2561_DATA01(2));	--16bit

chScale0<=chScale_TS(Tint);	--16bit
--			X16								X1
chScale1<=chScale0&"0000" when iGain=0 else "0000"&chScale0;	--20bit
chScale<=conv_integer(chScale1);	--20bit

channe0<=conv_integer(CONV_STD_LOGIC_VECTOR(CH0*chScale,36)(35 downto 10));	--26bit (ch0*chScale)/2^10
channe1<=CONV_STD_LOGIC_VECTOR(CH1*chScale,36)(35 downto 10);				--26bit  (ch1*chScale)/2^10
							--RATIO_SCALE9+1
ratio1<=conv_integer(channe1&"0000000000")/channe0 when channe0/=0 else 0;	--12bit (channe1*2^10)/channe0
ratio<=CONV_STD_LOGIC_VECTOR(ratio1+1,13)(12 downto 1);						--12bit (ratio1+1)/2

--iType:0
KTC<=KT_T_FN_CL when iType=0 else KT_CS;--12bit
BTC<=BT_T_FN_CL when iType=0 else BT_CS;--12bit
MTC<=MT_T_FN_CL when iType=0 else MT_CS;--12bit
BM<=0 when ratio>=0 and ratio<=KTC(0) else
	1 when ratio<=KTC(1) else
	2 when ratio<=KTC(2) else
	3 when ratio<=KTC(3) else
	4 when ratio<=KTC(4) else
	5 when ratio<=KTC(5) else
	6 when ratio<=KTC(6) else
	7 ;

tempb<=channe0*conv_integer(BTC(BM));				--32bit channe0*b
tempm<=conv_integer(channe1)*conv_integer(MTC(BM));	--32bit channe1*m
temp0<=0 when tempb<tempm else tempb-tempm;			--32bit

--將小數第2位進位到小數第1位round
temp<=temp0*10+8192;	--2^13  --LUX_SCALE-1=13
--取到小數1位
LUXS<=conv_integer(CONV_STD_LOGIC_VECTOR(temp,33)(32 downto 14));	--19bit /2^14
--去小數
LUXSx<=LUXS/10;

--決定小數點位置 (TSL2561 LUX測值最高約3千多LUX)
LUXDP<=1 when LUXS<10000 else 5;

--顯示值轉換
--	   xxx.x				  xxxx
LUXS1<=LUXS when LUXDP=1 else LUXSx;

--可能有小數點
LUXS3<=LUXS1 mod 100;
LUX(0)<=LUXS3 mod 10;	--小數位
LUX(1)<=LUXS3/10;		--個位

LUXS2<=LUXS1/100;
LUX(2)<=LUXS2 mod 10;	--十位
LUX(3)<=LUXS2/10;		--百位

--無小數點
LUXSx2<=LUXSx mod 100;
LUX(4)<=LUXSx2 mod 10;	--個位
LUX(5)<=LUXSx2/10;		--十位

LUXSx1<=LUXSx/100;
LUX(6)<=LUXSx1 mod 10;	--百位
LUX(7)<=LUXSx1/10;		--千位

--=====================================================================================
--SD178BMI2C--------------------------------------
--不同語音表所有計時皆由driver負責,使用者更方便
--增加語音表執行完,可選擇是否延遲一段時間後才結束
--SD178BMI2C_P_end_t_onoff='1'是'0'否啟動終止延遲計時
--SD178BMI2C_P_end_t_set:0~32767 終止延遲計時次數(1:約1.004ms)
--================================================
--00 00 xx --硬體reset
--00 01 xx --nop 立即回應結束
--01 00 xx --由睡眠省電模式中喚醒
--立即指令:
--以下2017  V1 版
--01 80 xx --清除SD178B buffer內的所有碼,停止正在執行的動作:轉成 "硬體reset" 操作(此版本80不會當機)
--01 81 xx --音量增1單位(+0.5dB)
--01 82 xx --音量減1單位(-0.5dB)

--以下2019 02 12 V2.2 版適用(此版本80會當機，是此模組本身的問題，越改越糟)
--01 80 xx --清除SD178B buffer內的所有碼,停止正在執行的動作,音量等已執行的設定不變:轉成 "硬體reset" 操作
--01 81 xx --音量增1單位(+0.5dB)
--01 82 xx --音量減1單位(-0.5dB)
--新增8F xx 2byte 指令
--02 8F 00 --Pause暫停
--02 8F 01 --Resume取消暫停
--02 8F 02 --Skip 提前結束正執行的87H或88H指令，跳至下一指令
--02 8F 03 --Soft Reset 重新開機
--================================================

SD178BMI2C_CLK<=FD(8);	--I2C時脈
SD178BMI2C_DATAin<=SD178BMI2C_sound(SD178BMI2C_IL+1);
SD178BMI2C_D_W_R_N<=conv_integer(SD178BMI2C_sound(0));
SD178BMI2C_P:process(FD(8))
variable V1orV2:integer range 0 to 7:=2;--如使用V1版設1(80原功能)(請不要下V2新指令)，如使用V2版設2(80轉成 "硬體reset" 操作)
variable SD178BMI2C_mO0_1,t_start:std_logic;
variable t,end_delayt:integer range 0 to 20000;
variable t2:integer range 0 to 15;
variable end_t_start,SD178BMI2C_P_end_t_onoff_s:std_logic;
variable t3:integer range 0 to 100;
begin
	if 	SD178BMI2CP_reset='0' then
		SD178BMI2CP_ok<='0';			--完成指標
		SD178BMI2C_RESET<='0';			--sd178BMI2C2wdriver1重置
		SD178BMI2C_reWR<='0';			--繼續
		SD178BMI2C_RW<=SD178BMI2C_RWs;	--0write:1:read
		SD178BMI2C_IL<=0;
		SD178BMI2Co_reset<=SD178BMI2CP_reseton;	--硬體reset off or on
		--配合不同需求必要性延遲設定
		t_start:='0';
		t2:=11;		--reset time
		--選擇性延遲設定
		end_t_start:='0';										--off啟動終止延遲計時
		SD178BMI2C_P_end_t_onoff_s:=SD178BMI2C_P_end_t_onoff;	--是否啟動終止延遲計時
		end_delayt:=SD178BMI2C_P_end_t_set;						--終止延遲計時次數(1:約1.004ms)
		t3:=98;													--delay 0.001004s

	elsif rising_edge(FD(8)) then
		if SD178BMI2CP_ok='0' then
			if SD178BMI2C_IL<conv_integer(SD178BMI2C_sound(0)) then	--send data
				if SD178BMI2C_reWR='1' then
					SD178BMI2C_reWR<='0';		--page作業:繼續
				elsif SD178BMI2C_RESET='0' then
					SD178BMI2C_RESET<='1';		--啟動sd178BMI2C2wdriver1
				elsif SD178BMI2C_ok='1' or SD178BMI2C_D_W_R_Nok='1' then		--完成 or --下一筆作業通知
					if SD178BMI2C_RW='1' then
						SD178BMI2C_DATA0_4(SD178BMI2C_IL)<=SD178BMI2C_DATAout;	--輸出資料
					end if;
					SD178BMI2C_IL<=SD178BMI2C_IL+1;			--下一筆
					SD178BMI2C_reWR<=SD178BMI2C_D_W_R_Nok;	--page作業通知
				end if;

			elsif end_t_start='1' then--啟動終止計時延遲後結束
				t3:=t3-1;
				if end_delayt=0 then
					SD178BMI2CP_ok<='1';	--完成指標
				elsif t3=0 then
					t3:=98;--delay 0.001004s
					end_delayt:=end_delayt-1;
				end if;

			elsif t_start='1' then--啟動計時延遲後結束
				t:=t-1;
				if t=0 then
					end_t_start:=SD178BMI2C_P_end_t_onoff_s;		--是否啟動終止計時延遲後結束
					SD178BMI2CP_ok<=not SD178BMI2C_P_end_t_onoff_s;	--是否完成指標
				end if;

			else
				if SD178BMI2Co_reset='0' or t2=0 then
					if t2/=0 then
						t2:=t2-1;
					else
						SD178BMI2Co_reset<='1';		--硬體reset off
						t_start:=SD178BMI2Ci_MO0;	--啟動計時延遲後結束
					end if;

				elsif SD178BMI2C_sound(0)>0 then
					if SD178BMI2C_sound(0)>3 then	--X"8A",X"06",X"8A",X"07" -->等待播音結束:等待軟體結束:不做硬體reset
						if SD178BMI2C_sound(SD178BMI2C_IL-1)=X"8A" and SD178BMI2C_sound(SD178BMI2C_IL)(0)='1' and
						   SD178BMI2C_sound(SD178BMI2C_IL-3)=X"8A" and SD178BMI2C_sound(SD178BMI2C_IL-2)(0)='0'then--等待播音結束:等待軟體結束:不做硬體reset

							SD178BMI2CP_ok<=SD178BMI2C_mO0_1 and SD178BMI2Ci_MO0 and not SD178BMI2C_P_end_t_onoff_s;--結束
							end_t_start:=SD178BMI2C_mO0_1 and SD178BMI2Ci_MO0 and SD178BMI2C_P_end_t_onoff_s;--啟動終止計時延遲後結束
															  --X"8A",X"06" -->等待播音結束:--執行硬體reset on
						elsif SD178BMI2C_sound(SD178BMI2C_IL-1)=X"8A" and SD178BMI2C_sound(SD178BMI2C_IL)(0)='0' then--等待播音結束:--執行硬體reset on
							SD178BMI2Co_reset<=SD178BMI2Ci_MO0;--等待硬體reset on --delay 30.72ms
						else
							end_t_start:=SD178BMI2C_P_end_t_onoff_s;		--是否啟動終止計時延遲後結束
							SD178BMI2CP_ok<=not SD178BMI2C_P_end_t_onoff_s;	--是否啟動終止計時延遲後結束(播音時間自行控制)
						end if;

					elsif SD178BMI2C_sound(0)>1 then
						if SD178BMI2C_sound(SD178BMI2C_IL-1)=X"8A" and SD178BMI2C_sound(SD178BMI2C_IL)(0)='0' then--等待播音結束:--執行硬體reset on
							SD178BMI2Co_reset<=SD178BMI2Ci_MO0;--等待硬體reset on --delay 30.72ms
						--2019 02 12 V2 版 8F xx(0,1,2,3)立即指令 delay 30.72ms
						elsif SD178BMI2C_sound(SD178BMI2C_IL-1)=X"8F" and SD178BMI2C_sound(SD178BMI2C_IL)<4 then--2byte 立即指令
							if SD178BMI2C_sound(SD178BMI2C_IL)=3 then
								t:=17350;
							else
								t:=10;
							end if;							
							t_start:='1';	--啟動計時延遲後結束
						else
							end_t_start:=SD178BMI2C_P_end_t_onoff_s;		--是否啟動終止計時延遲後結束
							SD178BMI2CP_ok<=not SD178BMI2C_P_end_t_onoff_s;	--是否完成指標
						end if;

					else	--1byte 00(喚醒),(立即指令:80,81,82):delay 
						
						if SD178BMI2C_sound(1)=X"00" or SD178BMI2C_sound(1)=X"80" then --00(喚醒)、V2立即指令:80 轉成 "硬體reset" 操作
							if V1orV2=1 then
								--V1
								t:=10;
								t_start:='1';	--啟動計時延遲後結束
							else 
								--V2
								t:=20000;--delay 0.2048s
								SD178BMI2Co_reset<='0';	--硬體reset on
							end if;
							
						else
							t:=450;
							t_start:='1';		--啟動計時延遲後結束
						end if;
					end if;

				else
					if SD178BMI2C_sound(1)=0 then
						t:=20000;--delay 0.2048s
						SD178BMI2Co_reset<='0';	--硬體reset on
					else
						SD178BMI2CP_ok<='1'; --nop 立即回應結束
					end if;					
				end if;
			end if;
		end if;
	end if;

	if SD178BMI2Ci_MO0='0' then	--捕捉SD178BMI2Ci_MO0
		SD178BMI2C_mO0_1:='1';
	elsif rising_edge(FD(8)) then
		if SD178BMI2CP_reset='0' then
			SD178BMI2C_mO0_1:='0';
		end if;
	end if;
end process SD178BMI2C_P;

--=====================================================================================
--聲音輸出通道選擇
--HP_R-HP_L及SPK_RN-SPK_LN(可以全關掉)通用
--全off後,喇叭仍會有聲音,可再由音量指令調為靜音,使喇叭不再有音響
--       off                       01:L,10:R,11:RL
--Sound8B<=X"01" when M776="00" else "000001"&M776;--有的音箱放大器可能會有問題
--Sound8B<=X"08" when M776="00" else "000001"&M776;--有的音箱放大器可能會有問題

--HP_R-HP_L		:100-LR:靠靜音關閉 :101-L,110-R,111-LR
--SPK_RN-SPK_LN :100-xx(可以全關掉):101-L,110-R,111-LR
--Sound8B<="000001"&M776;--ok

--SPK_RN-SPK_LN專用
--Sound8B<="000010"&M776;--8:off(可以全關掉),9:L,A:R,B:RL

-- ---------------------------------------
M710<=M70s(1)(2)&M70s(0)(2);--功能選擇
M776<=M70s(3)(2)&M70s(2)(2);--聲道選擇
SW_CLK<=FD(18);	--防彈跳操作速率
process(SW_CLK)	--防彈跳
begin
	--M4..0防彈跳
	for i in 0 to 7 loop
		If M7_0(i)=M70s(i)(2) then
			M70s(i)<=M70s(i)(2)&"00";
		elsif rising_edge(SW_CLK) then
			M70s(i)<=M70s(i)+1;
		end if;
	end loop;
end process;

-- --------------------------
--除頻器
Freq_Div:process(SCLK)
begin
	if S_RESET='0' then
		FD<=(others=>'0');
	elsif rising_edge(SCLK) then
		FD<=FD+1;	--除頻器
	end if;
end process Freq_Div;

-- ----------------------------
end YHGL;