library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tsl_test is
	port (
		
	);
end tsl_test;

architecture arch of tsl_test is
	
begin
	
end arch;