library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dht is
	port (
		-- dht
		dht_data : inout std_logic;
		-- system
		clk : in std_logic;
		rst : in std_logic;
		-- user logic
		temp : out integer range 0 to 50;
		hum : out integer range 0 to 80
	);
end dht;

architecture arch of dht is
	
begin
	-- TODO complete this
end arch;